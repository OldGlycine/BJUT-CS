module scanner(clk, I_ROW, I_COL, clk_1hz);
	input clk,clk_1hz;
	output reg [15:0] I_ROW = 16'b0;
	output reg [3:0] I_COL = 4'b0;
	reg [3:0] counter;

	always@(posedge clk)
		if (I_COL < 16)
			I_COL <= I_COL + 1;
		else
			I_COL <= 4'b0;
	
	always@(posedge clk_1hz)
		if (counter < 6)
			counter <= counter + 1;
		else
			counter <= 0;
			
	
	always@(I_COL, counter)
		case(counter)
		0:
			case(I_COL)
				0:I_ROW = 16'b0000_0000_0000_0000;
				1:I_ROW = 16'b0000_0000_0000_0100;
				2:I_ROW = 16'b0011_1111_0000_0100;
				3:I_ROW = 16'b0000_0000_1000_0100;
				4:I_ROW = 16'b0000_0000_1111_0100;
				5:I_ROW = 16'b0000_1110_1101_0100;
				6:I_ROW = 16'b0000_1010_1101_0100;
				7:I_ROW = 16'b0000_1010_1101_0100;
				8:I_ROW = 16'b0000_1010_1101_0111;
				9:I_ROW = 16'b0000_1010_1101_0110;
				10:I_ROW = 16'b0000_1010_1101_0100;
				11:I_ROW = 16'b0000_1110_1101_0100;
				12:I_ROW = 16'b0010_0000_1111_0100;
				13:I_ROW = 16'b0010_0000_1000_0100;
				14:I_ROW = 16'b0010_0000_1000_0100;
				15:I_ROW = 16'b0001_1111_0000_0100;
				default:I_ROW = 16'b0;
			endcase
		1:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0010000000000000;
				3:I_ROW = 16'b0010000000100000;
				4:I_ROW = 16'b0010000100100000;
				5:I_ROW = 16'b0010111000100000;
				6:I_ROW = 16'b0010000000100100;
				7:I_ROW = 16'b0010000000101000;
				8:I_ROW = 16'b0011000000100000;
				9:I_ROW = 16'b0010110000100000;
				10:I_ROW = 16'b0010001110100000;
				11:I_ROW = 16'b0010000000100000;
				12:I_ROW = 16'b0010000000000000;
				13:I_ROW = 16'b0000000000000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		2:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000000000000;
				3:I_ROW = 16'b0000001000100000;
				4:I_ROW = 16'b0010001000100000;
				5:I_ROW = 16'b0011111111111100;
				6:I_ROW = 16'b0000000100100000;
				7:I_ROW = 16'b0000100000100000;
				8:I_ROW = 16'b0010010010001000;
				9:I_ROW = 16'b0001001111001000;
				10:I_ROW = 16'b0000110010101000;
				11:I_ROW = 16'b0010001110011000;
				12:I_ROW = 16'b0010000010001000;
				13:I_ROW = 16'b0001111110000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		3:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000010000001000;
				3:I_ROW = 16'b0000001000001000;
				4:I_ROW = 16'b0000000100001000;
				5:I_ROW = 16'b0011111111001000;
				6:I_ROW = 16'b0001000010111000;
				7:I_ROW = 16'b0001000010001000;
				8:I_ROW = 16'b0001000010001000;
				9:I_ROW = 16'b0001000010001000;
				10:I_ROW = 16'b0001000010001000;
				11:I_ROW = 16'b0011111110001000;
				12:I_ROW = 16'b0000000000001000;
				13:I_ROW = 16'b0000000000000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		4:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000000000000;
				3:I_ROW = 16'b0010010000000000;
				4:I_ROW = 16'b0010010101111100;
				5:I_ROW = 16'b0001010101010100;
				6:I_ROW = 16'b0001010101010100;
				7:I_ROW = 16'b0000110101010100;
				8:I_ROW = 16'b0000011101010100;
				9:I_ROW = 16'b0000110101010100;
				10:I_ROW = 16'b0001010101010100;
				11:I_ROW = 16'b0001010101010100;
				12:I_ROW = 16'b0010010101111100;
				13:I_ROW = 16'b0010010000000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		5:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000000000000;
				3:I_ROW = 16'b0011111111111000;
				4:I_ROW = 16'b0000100000001000;
				5:I_ROW = 16'b0000100011001000;
				6:I_ROW = 16'b0000011100111000;
				7:I_ROW = 16'b0000000000000000;
				8:I_ROW = 16'b0011111111111000;
				9:I_ROW = 16'b0001000010001000;
				10:I_ROW = 16'b0001000010001000;
				11:I_ROW = 16'b0001000010001000;
				12:I_ROW = 16'b0001000010001000;
				13:I_ROW = 16'b0011111111111000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
			default:I_ROW = 16'b0;
		endcase
endmodule