library verilog;
use verilog.vl_types.all;
entity f_c_vlg_vec_tst is
end f_c_vlg_vec_tst;
