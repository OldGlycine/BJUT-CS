library verilog;
use verilog.vl_types.all;
entity flowing_water_light_vlg_vec_tst is
end flowing_water_light_vlg_vec_tst;
