module scanner(clk, I_ROW, I_COL, clk_1hz, stop, left);
	input clk,clk_1hz, stop, left;
	output reg [15:0] I_ROW = 16'b0;
	output reg [3:0] I_COL = 4'b0;
	reg [3:0] counter;

	always@(posedge clk)
		if (I_COL < 16)
			I_COL <= I_COL + 1;
		else
			I_COL <= 4'b0;
	
	always@(posedge clk_1hz)
		if (counter < 2)
			counter <= counter + 1;
		else
			counter <= 0;
			
	
	always@(I_COL, counter)
	if(!stop)
		if(left)
		case(counter)
		0:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000100;
				2:I_ROW = 16'b0000000000001110;
				3:I_ROW = 16'b0000010010010101;
				4:I_ROW = 16'b0000001001000100;
				5:I_ROW = 16'b1111111100100100;
				6:I_ROW = 16'b0000000010010100;
				7:I_ROW = 16'b0000000100000100;
				8:I_ROW = 16'b0000000100100100;
				9:I_ROW = 16'b1000000100100100;
				10:I_ROW = 16'b1000000100100100;
				11:I_ROW = 16'b1111111100100100;
				12:I_ROW = 16'b0000000100100100;
				13:I_ROW = 16'b0000000100000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		1:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000000000000;
				3:I_ROW = 16'b0000010010000000;
				4:I_ROW = 16'b0000001001000000;
				5:I_ROW = 16'b1111111100100000;
				6:I_ROW = 16'b0000000010010000;
				7:I_ROW = 16'b0000000100000000;
				8:I_ROW = 16'b0000000100100000;
				9:I_ROW = 16'b1000000100100000;
				10:I_ROW = 16'b1000000100100000;
				11:I_ROW = 16'b1111111100100000;
				12:I_ROW = 16'b0000000100100000;
				13:I_ROW = 16'b0000000100000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		default:I_ROW = 16'b0;
		endcase
		
		else
		case(counter)
		0:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000000000000;
				3:I_ROW = 16'b0000010010000000;
				4:I_ROW = 16'b0000001001000000;
				5:I_ROW = 16'b1111111100100000;
				6:I_ROW = 16'b0000000010010000;
				7:I_ROW = 16'b0000000100000000;
				8:I_ROW = 16'b0000000100100000;
				9:I_ROW = 16'b1000000100100000;
				10:I_ROW = 16'b1000000100100000;
				11:I_ROW = 16'b1111111100100000;
				12:I_ROW = 16'b0000000100100000;
				13:I_ROW = 16'b0000000100000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		1:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000000000000;
				3:I_ROW = 16'b0000010010000000;
				4:I_ROW = 16'b0000001001000000;
				5:I_ROW = 16'b1111111100100000;
				6:I_ROW = 16'b0000000010010000;
				7:I_ROW = 16'b0000000100000000;
				8:I_ROW = 16'b0000000100100000;
				9:I_ROW = 16'b1000000100100000;
				10:I_ROW = 16'b1000000100100000;
				11:I_ROW = 16'b1111111100100000;
				12:I_ROW = 16'b0000000100100000;
				13:I_ROW = 16'b0000000100000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		default:I_ROW = 16'b0;
		endcase
	else
		case(counter)
		0:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000010000000;
				3:I_ROW = 16'b0000000001000000;
				4:I_ROW = 16'b0011111111110000;
				5:I_ROW = 16'b0000000000001100;
				6:I_ROW = 16'b0000011000001000;
				7:I_ROW = 16'b0000101011101000;
				8:I_ROW = 16'b0010101010101000;
				9:I_ROW = 16'b0011101010101100;
				10:I_ROW = 16'b0000101010101000;
				11:I_ROW = 16'b0000101011101000;
				12:I_ROW = 16'b0000011000001000;
				13:I_ROW = 16'b0000000000000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		1:
			case(I_COL)
				0:I_ROW = 16'b0000000000000000;
				1:I_ROW = 16'b0000000000000000;
				2:I_ROW = 16'b0000000010000000;
				3:I_ROW = 16'b0000000001000000;
				4:I_ROW = 16'b0011111111110000;
				5:I_ROW = 16'b0000000000001100;
				6:I_ROW = 16'b0000011000001000;
				7:I_ROW = 16'b0000101011101000;
				8:I_ROW = 16'b0010101010101000;
				9:I_ROW = 16'b0011101010101100;
				10:I_ROW = 16'b0000101010101000;
				11:I_ROW = 16'b0000101011101000;
				12:I_ROW = 16'b0000011000001000;
				13:I_ROW = 16'b0000000000000000;
				14:I_ROW = 16'b0000000000000000;
				15:I_ROW = 16'b0000000000000000;
				default:I_ROW = 16'b0;
			endcase
		default:I_ROW = 16'b0;
		endcase
endmodule