library verilog;
use verilog.vl_types.all;
entity ext_tb is
end ext_tb;
