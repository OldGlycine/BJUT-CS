library verilog;
use verilog.vl_types.all;
entity test_mips is
end test_mips;
