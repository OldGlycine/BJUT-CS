library verilog;
use verilog.vl_types.all;
entity D_latch_vlg_vec_tst is
end D_latch_vlg_vec_tst;
