library verilog;
use verilog.vl_types.all;
entity im_tb is
end im_tb;
