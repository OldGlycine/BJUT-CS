library verilog;
use verilog.vl_types.all;
entity tstage_gate_vlg_vec_tst is
end tstage_gate_vlg_vec_tst;
