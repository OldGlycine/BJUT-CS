`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RYuoasXcTxqZl4OypfcV41Dwu7SB3dkHbS3Cg0LFsj1QL3FtzeIRLNOj7siwa8I8T2D4oIY5scPT
OIYHJqI0EA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c4RquQwHuC97o/rjIkwSApk/EDWuNTy6utZSdvrJqtGl8bh5FWGoojLTXZnMdZr7mYJTQp9fQHpp
HR1p28pRc2JEaj81rtfPyEJdSxz1D+830VGv1nxuRebLwPIiesN68abmxoPbFChRpgibQbJOYBIr
ep70Hj4GOkFunX6k/oY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
r9X4FEpeftZaomzB7fpgYpps40t6c6MJRatNxnTXgNtJi0/qcV2fBXUrQ3thFBnFDzIglq3o1gQP
3AqRJJM68C6x2Da7CHIQkS9VGFDKy+qbhYW6QunksTEzZ3pMNDNhIJCJVKaPu/SdrtiY9kSqeK65
F9vIOmhQusKrhF/n2O25zp+ueG0/q6o7rVrYb+yIh2D4Y7DfgEkC1HSLzJwY13Xdkwvdu+SH8NPu
jU43IK8CpDJ6Thzrp8ek94KdHdhksWOtuG++IxSE+t+0/ZGO1bE3WeedfH/wpU6zVxDf6N8/QDoM
wsaaqk315/NY1QG/ahD+U5hOlBWTAIwXd7u/mQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oMKNfXyneL4p/ztU77XWHi3an+1tg4h1hSFrpp60j3DscSF7r5de0GfsSY6r49E0k95gZKMl64AH
1m9U1HQChoj2WLJMUwPqAOlLniOdLUF4J1znn5xYWdO340adDpDHMEPn8F3RFqLPwQLxRtcP60fS
KlL1e7Gt0EZG5WFXeUEE0G7O/TlLJRgZHs88DM53qWPH6dRe1UHF7e/29l505cEN9BKz0HhMUoMR
XEJwN1/szL0xqs7bEq2OcS8gr0SVfMKSw34u4kJ59tuRI43bCYs6xwolLag8bF8GA4ggX/03LE1X
NhDhKnjFNk4pksB+DejQcoGXMPx+RyILpLohIA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VzpnFpMOj1x8A+QYv8fgXtvioP+QqCbRn3LqvgMI3LHpbFdc5UQ4/K0cgdlFbwSGet/Fkt7Z3QPK
1UuGcBohDgvNj3XBFE3XfR4dwy0gKq/vVHD4gXtRf5UHeDtwSHg6c6ii0X0Iv2coI5bV+iwh8MxZ
eKW0i6yO94O/UsseyRmJDg7zumPWsJyNB2+Se17N2rLp1ZZ+Fpoqrl161TUEtQntfHUxeg1a0emb
VXJbSeuLk93zciARyc5XNwp2F/lWO+dAOHIVhi2wbbg+CxTlxnLgYBbE2KnvHFFNXUhKSLmp+DDR
+y712hQR6oTVXueG/kc1sLiU14FRC41zaSIKkA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T2vtWi4yVyuAMDCgRlcOYSDYeCQ745ugoL5XAxPRQ55x0orQCShZ475xlcqQXN/z0iAOCRYE+9rp
5GM0ga6dsiYsXaqtwV9D05pheB1vJPHM0GsjPe0SVh/zNp9DiGmCJwuvzGYWxS9OfdQUolK2It/W
eTC/M1G5P28HiZ6mo2E=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VLywuJoPfY6IoEMvT3Hu2J4GsnExnr9ttNgiROyfi7daULbXwsrsvLjPhOp35sgcsp5sYKO417QX
qToj+PVFzTjVcJdVlwS1OquA7pG5xpG0QTFiDCHxmzvRws9XHzrC3lns91RdtQ+oK5da9LqF17su
3zrGQLgkajZEO3sAdOo+c3Hm8hCtKL7Fpw9+D9GBMkyFPL0XAME93srKKEg2dnpBP9wiqAAtz290
e3NYFI+kfc8JdO86lrneDXywb7qei+NYBvlo1CabsNeOJE2IIB3+/MIpa1Tm8UL3/EPX0F/0h0UT
lqHnjXlJITkLWt0Dsommkj+4VdxJKEc6AwZz9Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
Sutg9JR0Di6oMZx1GI7Lwf25txsLlZUH3KP/FXGerFQGsWU/gGC2aD/es211AyqmWOArZ4/mVmaR
X5FWnyPWNpyVm5DRrjdDVhXzFdPdzVOftM029Pusw4z3vgXj/gJWvs+3yN/1pAZM2TqX5/WYEhuB
p0gwfnS+NSy77pJQeWZZXXb+PVwnTJ56nfxOx/yA46+JCgoxaR3yx+4l0rp1wDDIVKqNrnZ/6O2E
g1Ph1cP49B9Xg/XFeI0rEFWDHx/3mISCod2q0s5DQoXA70wHslRp1Ho/ICehzdEoNK6eislEmpNZ
r9jnPAhw7UdV127c5w0ltlj9lamhIFaiphsJuci4GMzDB4jGfwKieC5Q/De3F1BgTHYwOuimTkhr
f5jKQth0ulgz3GMAKwyI0nTxiWb91TajmoPIE46lSRLIfUvQExFDvN0n4GNqAeeOyRKu428kqab6
v4lrZjipYo9DPmKojACwU3n8ruQXkl9YzIn5AOA3YBH+AOLeLRSL3dbDDYRiGj0q+xYN6RrUneLb
C8BoJLG3bqJGcTrPhtAIAnmjbSh6x6Rkb2bFoT3OwfawJBS105l6rOnWL3CgmBKnkuMQJzjt1lgj
Djaps61aIyXp6lenHAoPVWYDOBGxbsjR00OiTc3HUx4og3m1iTbQGqf2ATzLFL+5BhO1OwvlBLqV
k2ImpA7eAyvnk78quyZKTpTtI6nlX3TxgSQxqWu30a1CZ0A3I4su56l/aua/gO5u/Ku5V0O4lbqz
D+GVU8CSRSsWmNc/LhJRYFBSARW75b/t7iJKqkHcoqkTwNFL6uSfk++NzY56pFrizPLRpwpH5DGb
4CdVZF5mcy9Pi03ez2SNRP88INbEo+/UxoVUJQ8H/tUoKV3zBPDVvHzW9XqE5xUgnij7uh/TzYaj
bE4q/GgJuiTRBJGnbcQVmqVioJgzqTUcdQR4lmJjuTlgLViTgvivv1rjaFQHrzB7KJVcik+q7Rub
lqiBIxjgtg8wfsDEUt6A9kGXo0/BTNzbWNnATOd4XAQfiYEyOJS/YY0T63wdandMKLEQnkYpUSYJ
aWWeEdV45ijUuFCBGxHIOCHopn2WdOpdt/ao/0n21sdaUnhBcMLaOAgYdJDfP1rp48g8fI7w9dB3
erBZ2xzxXq5h6WfiYBx6tOqVgCtXBwgnpv+0Abk0oLRiFmTn2pjXz7xRIB+5J0+GLbRcJNYGFlSS
t/eXcF8iI55pGdh/USHvbFMN5tsrtEV2d/kiTXenb/7YN4ElPnhAQkc+4jB8PZvi+GRek7S5fijk
QCH3Qfz9gyPCsR8YiU4bhmD7BnFHqcgIrnwL6lHJOha7UfAClWTSgoE+qe5lPkdCytwgRdFblwPt
DO28x+/KhuSp8Svyu6UmthjM6ZzHIVOeQyW0XbhBvik++JBHmg6rgY2RQWUw5FweScDw0ntUUgwa
h45D9cE5Dgz1KOSajYFJphrNSiiKrnfMddgBchkqTfmLekioCuQSfNCyKREXxg+U7JzqQ5L5MJyN
u09bhUjwUvPuM2r9xW3pdg5NPVwoGNBSgbw3nchRInj1X9BUvczLjve9DcWd3V5mh8SV6YYdXfKG
mfLYF0XIamwdTZ5p3tr/a+d0+Srsgr2/OkdY6Xm1UAxZda5aMvzvEtga14ttKJ1GOJWZICGV/vNY
4uF1Ydk7mYL3KdpvbDYG+IciHijBoGRxGihkhCFjgsx531Cvv9HqTVEf1yYWmEPAnD+d1ade9OXi
cCOI1DxolNkzvHy5SxTkO/xqJlrVZwh3PM0pqm+fBM+J6Xr/ZDyL/Bj9t/EkKl9t2cfDhqz1izvV
b9epAq7SyYYpMBOtat+DgNIHtMjuK8/5DPcGjhWFotpWZeBe6DYlABaHLaA/6B5n7B8L2ebtAskb
5B+SLAuoK585/kydVcWUXUUHwyfCqi8KT2vK2FGzPHtglHTK07QMl0KL0oETDp7CxjztH7flIoEU
a63/LFcb1S0uUMwa3nf576JwgW/AOfhs1E/zOnLG5Biqe1EJ2TyDss7SIlSIxWg7tr48OCBSc0/i
y/ei6bcAHYWEENAhwiaod0bDvBcVgW05W8dAZSSjMuAxhaxYe3YM+oadbzQCVFyYkXsmEyROIHdj
IW3o8XGt9U35wYjqGVeY/1rEWEk4aAvTjJdtyRc+eJsSM51JP/FBucmbHxyqWm5rKGFIiKl3nW9o
sY+QuLmvz1nu9mOhqyp03mlR1gG/aSEsBnH1ShYsGzzfbdKUVds/4XqVz8QEmuu5UKZ79VI/Vnzb
Pu+79bozZnaCORa5EeP60g7dFCc4CyfoagIny6u1cmdftaf+Di+Qc3OFoLypQEBz5v+0QPQ+CgDJ
O2CxUsS5ripMMqaoc62WBmi/fiJsRLz4BoIAX35NL2IAr3zjIXnK8LO1cyAfQO8RSoJ143fR7Y/M
thQszxbsFYE5GZXDbCTDLtgTDk7Wps2lQw91dAGS4/tlf4EUw5/exuakk3XfxcoeJPucwntZ1ygx
PxQUW6+J1Xr64K+t3yjMwmKF/lS4h9gjp5kvqu/fO+wF0LR1QtP6kDUmdWs4lehSVqcKJ6iooCDH
mXCWx00F7guGeoIykEFM1Weeg6q+LwTbL2IXWzLwzFRkLCxeGw+DHgfwYPAeq5gnxrgaW3Uz2gTH
DaF+VTLg2eGhR+pn2JM5ji1cAKHo+3bqReP/F7Ndz81nuhqwg/zuv2n2pDoA5pSogMHZIZ0ejYTb
Uj2ndROG1w/R3w3q0/EFWIcgytlVuiLYq7V84idqRGHKM5+Mg+/G+iU7LlusMIjJPXRxoFrmxZIq
Ni92tWBzxM2Ksvfp4eiaLVsBAE/bvHci2eykOUhFFZnnUOO2WpZOj7KUOTVwn/WI05iNxJZA9U0Z
MlnlJImPdiwhP+9IXJrLwBt228OwyPgOIEikUSUlgRnQ5L4bBvUYW48R59d+549RnoZ4H0E6CyKC
ysySuIk4K6QBuZVPMBHh1UyVZuZqd0w459rE5o8a9XW8ODAUFF2Je2t/GFMW3BAXqxlsyLrXZty4
AL27tdsRn20OWe3l4WcEAah9wroWCvAXXkH5ztXxB2c7ks8tocfjXo1jonUfZ8zVJjavL28MrSMB
LDe/r8sZUv5JsvUM6GDzwdMA4ugO0sjAI4bD9KSbpW2zW7kZ6FYBVCRFr1BvshmX6a62s+xXjmZn
Z+9m6Lv1m4Q/o5MgXWsTC1Orm7gMhsNUx6FoqjuM3Qh304zxjJCLByUdAZvb0OoMvgh7/EQ82/V8
YfnxFhhCxPID/Ht3YDCB9iDnRiwAl2IeDfADDNxtWRqxOUpvU15Jhntjvd3GLc94vqYZ0eO25A0s
mlgX9WlIQ02ZR0QXNYepg9eU3P/qvP6Oao2IEold8do1nhJ8a67WxW3+hnuow8aCjWcUgaLkGaSy
G/jjTHOrZmcBX9qcUVepkWa5lDWu7sEMUF+3Ub2r8OaEiUKsgUbh5Tx89m9szae+k8efeAecw5wI
UwWnUvQNFsq/zt0CG2FrmM8j8GK+M82kpJrhEHCaj8Jv8MApt4CRhVNUCm4DVJumXLq+3pWbbxW2
lY0gU2Q0S4ens8B/q4e86P9mC7VIKKO+pz1uRIQSculIexJINNP0rAMeHmcP2MzhroyzFYmKYhRn
vCzw6UwszG2PU+JrlXG33NG2Oeyi0ZClgAy0WeLi/uKdrvXmzLwDIG5SnQWTTuz+CROFfwsD7V2x
RIIqe+AWLZX033Z/ipmnC3GdDez1oU96BdclP176L+ilpPLxs30JQieyejHpkeBvwF0ua5GRjn8S
RvpEqnFImwzU83Q+yVvJRxsebQ0WUGUEgqPyz88NYCBE4ZOaLWlCjcZvWgrcj+BNYJKeG8kGJPSj
PMc7dqTExTJ84dZnwbePfwpdL+s6/w/BQm40o3RhJjUC4nVD1I1iLBhiJeOyllg5DJ45j5QB9s5i
kdkIlIJbCWenGzmNsPwGlBGVY4LmnSkLtVoVVWStNjVfAbiGCda/1InLbsUb7XzT61GbgN/0rJlg
yDPVcx6QSET8yA8MJ0YB0J8srJyMcy8oh5HGwFf5rFjaPvoz1J1k9lIM0i9rB1sR7UX0blnh3KGn
6pbRfGQR2xWQ4cIjbRW1V517kviIN+6EexZnEl0tMr+tJo/fjxQlJytKqBaO0pVfm+9uEjvxiFy2
drxFlTdSLnwqB/7jHdWg3Rv/I7956eKxia4+NMVj4oJIvgLrKrzqO/EF9nmdq/o9SeearxdomliJ
6Z0+lyDPXAPxyZHnnOeo8Ys0hXsKCIyCwvByWgF7MF8R+qvafxr7XegjNjv0BdvIEnCQr/MbaGVs
lA8os+bvr3A3tYSSrsR9adq6ipIMVGcwXeqtZ6WUAJZrB+YDyVja7LiAogT1coAA6a9ERF2+4NNP
56az9GP6s5cCgt7duvboGsO+3fcYvhqDb56mnLhY22FTD3DlpIuLcgr3+eFmfD+9aQKoq001Jl82
Vgt1AoaJ/uR0Lt6zc9ko5U0D4pVl5+Vr4M7UXOLH7AlR0iAg13kCZF2YkBnJBEydKl3nE26SvDx6
9BdrbCBCbptfwoxfP7yGp5aPM2KuPOp417D8a5DPgRfUNs0EE5lU8YdjcB/XblESLwyhvyvBn297
A2Poz9uesdAaDY2ztzQ3MPg4/jb0V5qP9ISt4GJYeihpHirMzCK/0UgA1T+gm3npiCz9SXXjqTKr
oyantnncvHtMbPOFqSq+DYxSfwDTCDaIUWyH4zSqtDBJg7t1oY+1ROhgqiFF/GEnwFS44eWU+zWp
MMeVkZjTT17l2yyG5S7xv0uyQauciB5mWUqSRQ6+uRS5H9B2ISOy0w2X44UTKbFXH5LEUcV3n+AI
xMbw4I4jz8AmdUmZ2sTm1MpGKnO0Hb8KoBEjPibD7SGWIlK9ZQZMpH7y5dgA8WtAG8GrgCMhn+mj
TPkFBFMUd8bZNdDpgZENyksiLdVcdddd7V2qjkyAhBQvvIGNsvu0fmuYhsYolRty4OtUYRgCczuB
UW7bghtJ/7VQNmJAT1+RMheOjIW/NM3da75laH/Yh9QDncE1p7KeSL3YFoTuBo34Nc3uNr7ilNiD
GZLMnQZBRo5VdnuxsDcyfD/Ix4VkvXDbMobInRU5fEl6gEy6zudr0UsgXVkos7y4EljV8HrlhHg1
R2LIm2CnOgCLaaMzXrqrPAhOWRRbwxx0bV2k1/5peWNZlFfChjhTUwz9gqZfygI8ZRObc+NBfpde
6S6XKdluu90/jkBdgKfpvb+NXz1fXdeSAtNEnLK7W2yJFT+92EvksRia1c8aIGNrTOQfBQ1X2Gna
MYXvcoGHiQ9drmj6xNTSlvYP5t7szuxtz1PMJJc+CgGRlJDrefhT+6H8h0tbtP2ZKoJ5ZN1PFNl6
/hJ+C9IVfQVQ4L5EPut3Yj64fM+UKBpeKz+ERniiC4zIAO6bq9JSAYSn3KmJG3Ovy3g5RJLpBHlz
n5qmmDhrf8UbYryDgaaWTHEjzdZHsiZ93Xot8JSoLe86jAOKPFPnlB3V7y8aGpYP8J7mRNhXehK6
OUDUWkoS4RidOxMfXpc8LqpNhbai2m4IKj6qeaNi5UH0HRp9uZ4mkf6uKxM72CV9wZvt7VsJ4wH3
Ean3PHBnLHwh3RP1+1hQ9i0dlp6sWQz7fGvLHQ5UQM1jZS7c4aSc+UAHXWMK2fJX88nJZ4S5TmSw
W2WQ2gjq0cKwSAfwCjisyQbageT8bl2Da8r9aDkiZ7LwfPqO0HZSolccPThO+BG7V3Et4BPW7j4o
rEA4FinCbBgEgn2rY7vM7wAPLoWMion9SiBdhovugu6vTwmmWZg01os99IqyCgym8QmNuG2GhUc6
Qgk0SlVC4I9097J2l/tNirVsYR+2xf/agqVd6iPA3jW7ypa2oHnQV76go0tlYLu+kcEXFrF2KQnC
XxrnjU+ldsEYeoJUMqSWu7bb+EcBHcX8Zgex8ObXbxRw5gtttJRBbPWbUh2U+0GbAu2qSQpSXFj3
Xx3q+oCCngN0jGuQ5RzjxFIX42VHOuCrbH85rqIPZRvNP2DNlfvbIAHwz5t2PtYC9ZcqoQxGAdS5
1rOD7XkSVIHbgFwmSc/EuYTRQSenQjvdbtWs3QC+0UNr7+zAFzOa9QQGI9joU29DZ/03U2qfimwR
jT9T29ldteZ4X5OtQyc7ZCfTdDGDmR8Wl2avsZBIl0XuDnZhRrLygCm/qjt6J2YHZB4bdDD4gW1V
hza5+H4m9FCfcq62eiV0gdCW85Ih3jBWaG2E4+YzIGBlGk81+nYjHSpXqctKEAXTt66y6p/FlNt0
Ya6wqFhdCR2XGU9dDdKDM9oinmzPQ5nyyYrmoH1yY0ZfECwim4OV9dQ6vaY6Ocy0GlFIQgCv+H1t
SnQLPjQohdo/wP81AuhhIs+edPZAqS/0lFeq04Ymx7J3JZ0QxhnXXnqqpum6C5HF71rXVSKFV6CV
zpdU5OlqKM1egxQTloqwrdaF5tm73XhJCBNAKtK+mh+R3vBEuyoqmLMYNfS9d9l16X3X7e6316XV
ZojA4m35ktu8PXyQFHdDDYBnEbRlziPqwrNP7Che/4GDoHdZALUvb1CHzDGlqc6jgIvMEFStCqwq
HEdbmNVXgZMKzKu6CAKIC5GuA6KsqCZNbicaHk1n01NlKhm5Pu1mSAFNQ7biRLoYs7zZctcqNP3s
LvIZFPD7SAzti2XSj4pBRsER7fXXYoWazO7JH6O6NEm1n64WjICoXwFD4qt84gtMh9RTs1A9APCP
jKmwFyKlH7BnHGGk2dvKRzQFJuliHmjfkuvttkEPGpbLUFGfeXah51tIIyQ8hzku7RklLFfoS4mW
yG4bIBuv3HaZR3tSnttkBXSDdFnAOsbX2+zvaJiGtkjRvotdmftAlUmstTxK7jtWV5GNpzPpP4+R
0OGQnROgBS4dFiE7HJgXG8ErDx9hRk94zk/SbyrC/p20iAkFAYBn0lO7mmCg9Q5JRKESYuRAAAYO
/AyfhZpWFHX1+FUF3chY100jbaVAl0b6tZiT9dJujJop8VOouAe/NbWScc8wp9yf0h5febHq/Ysf
ViXWHYMClpyPrd8EgLJlMIbprBVecvrkbq/iGGE6OT/tCRIJIFQch2+OstgrA+PX7k39arre/077
oHyfB9iADmh3lfzZf8RiD7O9ayWbC4df+M23y8ifci19qY+0sL5JF8SVuCvBCUoOQfi3I/dzFsxS
K2pSUcKm0SGGLM1aXEDykDVdHNyO+beQdNPMdX6R2kn80OBU5LVcw8keNFUfjzQQ1wIL9CtfHOqx
bm3QiMazFT8tOl+ebzqe5dD5Pnxxo1VUIqjAKd7NpYIL0xJ39YfNVyiLIijuf/ZDNdmlm0n++gtr
tnY0FQB/tRh+OVoFAgv9sqj+X/PDS06xsbRH50D0JJ9lhCBPccowY97YkPhn0c8vP+7s+ILKJfqP
oakNeADMI9/xwu0wHQFO3l+e2TB2CZHgc8u+AsXR6u9CrZSCyXN1FwXl+J2RPyJRL/eoNMAVpIuo
Zo6UpHxizeEiaBQYkJisuPXxbkKZAfSELtLFWLOair3RrkhaLi+HtmyCM4JOpK4V7799KxRpLJ3I
Wyh3gWyf1zEy5drvAEYp1wbhXM66hLPZCPVesJy1MbQvvHO8SN/8ROhdYFlcT4dEjvXurB9e2xJc
5PqNmjfi8CgK3hNyDTXGqSAQsZdE2HIuKRNJSlb3GOy6TJaC4aFFh7KsrR0joSKLxjLG2qIwNQEI
5qEBzJ/4Ni1oP+YY4ePP0h+oG9rdXu8tChC6utLqMoJNaB0VOZUSxB+kGeXywLYoH+LtKtk1udZS
+CjFCCctiOzzVLQS0tHYnTufTGPqpBbxpixyFkuJ7ZczraSGMn4VwSV1Q++7xIXA95dYu2SlVvnk
p8RpQ4kJXmnkqdYKmF04hxfYzm81kaTl0L1Cc7qM7H01Wi6TKXIJoXbUxge9jxYaUIowmEUjpQSY
DVdtzjTQzuNgjrpsxg/0Qma43CFfQ0SGT5tyRPeJ9jMcNmNb4zFZ5ubpwkyu2HpBpB139kZ4qqOI
ir6MZjEOs43xBCPaB2/IY5IioFjQj7cm262ikhiCLdQy2d9Wpf1fJLQL8wS+PzkszUBMdls0SVxN
ZgJkWb+81WVOljJ6QMZYGEa36DR4AC5RNOpFT8i4mAK64iH35PiVNDArJzZK/GlCYQ0HGLI2rVqg
wz/wyPP67VWcU30CxOp2t3WMBhkElOtk65pyMWBy4P9xRq6FlMAc9kJATy1i8ZnS9i1yuO8Mo6Tc
Y4VBaRuvo7TtwZxEAR3cyPkbUSJiEhEe6JGXxzkuJx4gfJEkRDkIAbw35HNnzvfLFSlW94L0WMAL
b1qOtmbf6iDn8nY3XjmneEXMtqG63YmCuxnby+39Vp57QEL6Xzzo4toKlAuU5nl+/CEqDfZKhPAg
v175gE0/+Eee+J2Qjjt6NHTRqlIbXK7cmcFJAbStFVCp862BTxHeTPs9urMAmawxiwAYa5GYZrLc
OezrsG6KdR5sGt5pbA1z6Cki0oWfV32xDoDVoi5cJzIuAQz6cgBZCQ4IplxhwPJpx8uzddRP9eYh
ZgFUSwhciQGzcqAyxJsWcCzHLBJCVRmyDP1pTvhv9SoRzHiLaMJlneLKsTmiguz++crLraitJNYR
lKvTrbytODoYhZV5ho9IVNKJb5ShIU3ct3rI+64JgFC+B0dh//m39csbiO0MtyE6w0sMZ/7ut8AT
kPIzYbbew2QuGkqriZ5TL7mxc3xHb5W0E1j4+FdCRAZoBPfZ9u+rFGhPl5wiRLgnwrUloVkZy3b4
XjQotZl4sIzo+jKR/DQ1ig4ke4mQaPhR77W8CXOyXkGpKFSpOivWWHoMuFj1saKKIE0ciFl/sI/C
d++/Y1e50vuCSF5YWKCwCxFHCKPExkj7d39gGP/wWpfrCY6oHqFBuUzl1S2J6zLa+HbSH5f7IyO4
IdOxLGMxoGLBnjG7UCrTwXsou01jtnr8X2jOnofJlaem3PcAkuZ39WW8uBx8AYkCj32BcoaOxILn
aS/usSFCgpPxD2X2PYDcLHus0i6VweVey1r5OinXQyRrxgCiIWgzFEyetQZpQD+CmvbvQjHkSnWt
BGqWyAB/6GPXhmNFPKVWTFjAXWd/vyLfryGO0kNkzlQ6t8kwZz0w6E7jm6GvDKQcDWvV3LzzYis0
RCBrWq7JeI8eR8NBgb/FvdUS2ddrSkdU6eMGe2hroiDiQUOWbXGfpHnYTHcYd0SCY9KHCKA68wr6
09WKjkfVKVwF1gemrkmh6ci+NLKndYVBIhyZNDUi0IXfDW3iWTCidwoAt7VkAuDMyy165snqrevx
WY79Zb5Hcj6FI1wtO3R1djlIBnj6anTQmu/oPvWScow17yA+jwmCj8zwu6ES915r/ZkeqkaQ93qp
f1FUrGuvifnNL3G8Qb9zBdJ5GLGGIQOx8aCrjmTJzM15fZqDvX/FbfN///meytIwAhpKsiUdzBWO
bmh8Qo8/W/pxt8pnu0GLcWFc70dNhJ7Q7kXak7BUJ71uMOwqlpppQeolyzyHgAIoPPdYBkYKfJMb
yOsmTV3628BFmZHbMzQahHVriSvNTA5GHTCMZIPZfjh5sRqd0MLmVwGrl7mXd7bvZgU23UtRd1xb
AXjrLro6LAULq57P6FdJobOPFJbaExuWoyHlT+HTtsBDSZRqO8CFTe1sOPhbUWbcx0gSoaJM8wK4
Y/Ubc2VSNQb6BiwqPJx2i83yGCmGeb4t30rwzg14qC/YZft5bn9sReHUrsPl24s5rClKIlkxjOSD
mOsF4pphz52/V+zj/ACBpWd25F0m2Br5IwtXx5RTEsO35q7TDHkKbWxZBOtCf5vfxZCkKHzJQICV
HL5+Lc4p/LRwck4LM/iZQqM9HfhWgzH3CtLCAghWGHU0p66mKFywNYgYPiwYiUv5rgQg7od9+Acr
jMf8FafnrwFCbOUWOF5+fC/qDbJC/bfx+W6rSucUSUP8UVhLFPck9WOxV/UwL0I+y4WZEmAmxpV0
FkVEZNtGlHKqL80GUGiZIdGEURsAq6IOgrCQ8xKTrS99PcY7I8TAbJgyPlLwpFgXNapCD3Eo6RRM
qYW+FX7s2sqnTH117VAh2ShMeok2F4GO4gjmXfWWASuVkUWcH1m5q0ZgPiMb//Ye28XN8j+iLeiH
rJoHcFBebRk/Qc0lmyJRxZdH+v+nlukfcG0fX3dOqX57nwMT14Z+UVVzSrEuiiuZM0z3UtqSE6Ov
sPN5ca3QdoZ/zq9/uVKegksR6iut/bGB/UMt637Kqxt26sJfGNEQwtxX83pgmGt62ObYPx4mF9Sb
hWz1PsC0Ffu8xNzKPlz6MP9vuMnjrpiu/aVIELqKfNl7avSEEtfCfirv65iH7+1DVVr0SCT6xAXr
3QCXF+bO89GYXThbQ1N/gvvBPAGehZBheNpn1WPfIa851/CPjClwrplpWPf1OgGgXrPC4el9BTqh
3W8WoGEruAJuJNNG4wMLgZIPTUXiAeQ2Qjm1Dob0NTvNQXapmyIW8IJwxXwuq0jyh71JxYgvlYqx
CznKPa59al/yajuZXkgrHm8x98C4jL9XFc9kkFacelvznlCOYrEyRKG7GJ2pin1X7QPTsMff38s4
nt/RRZvK2IP1WbwqHaZdLQpH7lYUiRefMcM2Nk2EnScLgVyb/t37dmW5bmUT9jCiJF30qkwuZ17e
tscp4MYoUCmcyRGOiKrw87RKUjrT32UWTj7X2tyR6GMMx4An19ZQJNfckyQQxQCJFo14M9SgjgxM
XYf6mi6pybr3RtubPjgY0d964nk+biHyEnkW2me8umfItAZNJ2duvHzHwyly3N3jZf5AJlI/xYLt
hYkjobmAyMxiojphR6fmAXNix0I3y4Gc+sRi5tzSnr3rGOFEdYsHbjNpoh86tl5E+TWDka1Iw8Of
syGXie8nKzo+g/OkdSAaESox9cu+frI54Cv9+wphS5ZGQvknAXd2sWjEi07KGExIAgsIZ+TjTOk5
UTX9rjvK6IQfvZdmzECwHpzcrP2Se9S73pdVf2B7Z6bSOr63dQOmafcrRzFya7YM31C0/7ZQS4UF
K5iosXN6aRpMtZt6f6muIcbNiQxvypIp39Bn1e1t78bnhYgXgK3TZxuIM4dFn3ySbHRUmInycdYO
pVpnTZQPVy1cYS2C2/uXznPAqGXUY4UWqpdD5QWGtIi1qyQAYVmpTlHRQpTrTZERYL7o6/nshnVb
96Dzk53JiyAr0K6tG+AdEZtTCzM6/BY9QnIl8fZtmMIFsb7pFfgSrOO9FkgxOnStygiegRI+605v
fWPfXUh1qiFV+WHRKJUbt+63YovWO2faSlClP9KLGxKBVLaVAuVJEkAGj1di2ZXI/1YoqsGMZBN7
e/9T13duY8fPRwc+LGkm4E2ikFTZIoeVjqRzxGMQpLxVVCpAIeiGqjSsM3PyUatI01ZDBm6y2IBq
McQgisBsJjwEF41qhfiosjcnwmR6PpGXQINM7Q4zgCTs89hWCD6ISoYss6JD2eoiTqPmkZvtGnjg
0vFKFCKw0iM0Nni3gWHEnrSZ5GjTL/wiN5N1jzGjxM8BjuubsQBGwdwMySrjwHr5UmJeZbbuwcKQ
QsdC6HZ211m5WF6Vk6z+TjWeSV1I/OPYiLDqApPHns33/AL5jr6Q7j6QZwv+qwoTLvtLyValxQHB
6FjQvLpS7oTX10yrEwbJyPkQFUikCChTGoyRupy/5xa6xk9uDggjIx+TTunmEpwZ4qHz9c2O/PBQ
HWyyW3PlKyV7JaB3x7g0LZY4tfLEtw+nOg14xkpLHZlaDcllxkPL5+/dfbTRuvDfs3OE9wunVQ9+
wYmt96Ac2CB32laVGxC1t1Ux5gDThjIsMD6yPBNH7unHm/mGraxbbITQdJyA1z3gQ2gWx1yCP0Hq
lXdbmZr+d2hJyUWwl93Wb4wMJQ93M98ZH8SuZW8XjJKQlg6fN1BR/dVgEEAPHehMY/7gb0eGkzgy
k4psdkLdkVUZMBfjGi+VtUMbSKRALtMTOSXHILkCcAZXzi0YTtfkQUa3KCehJsuX22SOnXP2GtJU
S9w0sC3Bngntx8/xqF1e/x1o+tpWeDO0tqEwmkM0ZyZIP7gcCQPsdqYt2ODzrL6vaoVGBNV5WyQC
CkhDAndEZCFSMp2xA4qsV81nt2HlQJF6Wem1taZSXMmYKUqU/FznwElgb3IMCpWusVgVGnt0aJyL
Hfbpuy5NZFLdLdktUCwY6MEv3tSOeDDufz4GhvU+9DJB8CVOaUlO+LrZMB36vxOwZQlJHORuYXAH
A7rpI2P+C33AXzoApzk3CRrMGLPZffcVX0N2WZjYNxr4lJW4l/VYUrV6wXANXRHD/Ujv8LCWpJjv
uAf2CBaqzkst3y415SOqeysi6VoYO+HDuIvpBWUDGm1E7B4lyZ/eHNQMK2wLKAy6qjVCblk8pEwC
OhkPEWuFox7dAmrupHHKKFkR3PewJ1ssQvcPljJN8yS3XZQcgle6TFynJBTNJEfktyBYISRNM6iY
EaOuABAte2Ql4wBiUJlPyO8T3MuY+7SyuEYNQbV/oMsDqnRvvYa8xQTB000Tj9YhD3uTct9vEada
4AsZyCWHY8U1DUVK1sr+862Rfx+8aOFfi6DtHONMKuIeRuIBGFz6tP2ylzyqdl/qHIY26z9LEhNG
CTaHXVSg/Nf/WfBkLN9HXxZwVXk8nCKlDm7YU5qhpN/EP2lktPQTjC38pedqqPsrCyRKeFdkHKrM
A77+i80qV2Gbn5R+D3ZaQF+vfUH/9rin9e8wHfXTOtKANl8WWjtmf4xySSa8c0/9XxQB85FL89Pq
sumrFxyzQH9f/6iVUedXPsj1jNbdmJMZ+ACsMbvRGeoeSLNl2WbGfh/nAxyr6dap7mpYLCaQzzVk
HU+pLOwSqeTvj8N/oG1gBYiJyl43JEaLHviTR8yTDQ1Vr6OAjNYf24AExsD4vqwPxc26u75Wr+7J
N4HFF5Hg3lJ8K+Osw7wxhQhGbVQUAUsb008u+kdHXSCI8xToM8SnFKltqxAVVHOyyHoA0p3FkV8c
1PfaSpsrD+dS0KoTEFcPr5T1Jx4aElVkWZdbQluKfxaH87VeqaXEmNaPo0IO7qv42IqW/MUlCNPi
uUIaCiayEmqDM3xxvGTyyT6Fb/glgEVNBlEwOzqNMzL/WWvljB01Q9bV8aI2DljJF/dBS4vS4PMU
t1J6uduYpvj+3/xkePOGn21tWc2s+OB9AM4m2y9XzFNfnQw+yjum21DvMks/7G4BLaHKkq8rN4J+
OfmGfbnWXo18YE6TaWPJpxbzLuB8nbzP4sa+GhMfsK17PQeWegYxi//yT2mw9TZzk9qF+kHKhSty
J3Gd9rIRmPH0WZLgAq0RAxoP485elH3yUNJXe9r9sGgNLB88fHJxjgLZ2WyWOZOvAf/cFZPey5UV
GO6ynfjCMXwfVs2cfQ5mEW1Ue0dmpu5OEZOaNiqJqJ1GWTzML0FQ1HfLZlF+pVqzVgxcn2rawNoR
MeAY5gdfXeja2gTZiWTRv/mC35zl8t4ciapU1rrlQ/N07wiYAmkgd/jLIeSvjWSLWRflt28Prz4q
8jhE4RxO3Tf2zLGRjnFqUy5zEbXw31BOdfRTlZTSD9kcjDspc7AE2aHwWTxpbaBdIiZ59TmdZA4f
6Wmvuo9VUHxmfxx2/9KP/X9Bd5GCfrdMmlX/QFvT1joMAJuurzApNbnBnfwwmmU70g8XYx7ltI0l
u4XP4641+uJJLN8cewo7uPOgbG4Oj6Bim70sVgTmJ3TkMSG6M9nWKCdcycJQjoZ5tigxkU7zftmy
O4M0IuHaj/VVnJUztjmzsMtKVlTjZcAIRzzGVWI1RXJfX+jQfn4CrEEFeJv4BX44feJJlfHbuKmZ
d9XbIifLY/dYuUk04tOVxgF7Fn48YHOz8MjNwbC/qmeRyMpDJswwU8PwKATcn1/5eCWERxROgH+R
nevxPt1NsILu7/fCL2TQ3rVCMTp8Is5h073MS7stT44CUVzk2bJbdcAyycUbBAXp7Xni9+H6coYq
hl8bVuC3Th8Y411cUG4inGz8FIKbrURMGhVrvwfTuaJGNKDKMH7Ugh8k2B78BZLwW4ePwD3ErJaz
VMdHYFLlEtCHZRwXl950hdZPJLRkSYSUdxwpHJ5itc3uu6OprZMDKDetDiNE+CvdT4Nbr/3aa8tM
+Y7GJsI5jWGsEdi7CMeAK1HYo82tPBm+nySmL4NteWmPuJwxs+LWWv/sCeBM9mQ+eGs5C/+X0H2C
2clX2637cnV0m6cdh0PZY9Vba8xGBvOg/v9btP7vkCP12QTAIwhr/M4tCo6jaNHt29rGmJpCAQgt
6dyyDscWF8hrlIT3MbtHUmIRK8AB7eBy0dsiq42V+KXSN8hIQl+aumUVP9L0/KqSdD4ZlG8PSDbR
JJqI73ZJ/ob+xALiePTtlx9PkM8sUQ2Jtl1bQUbOdJJTTS2yDwDmxAxnzJ+pvdZdB68T9exU2Afv
FK62CJ2l1gcTzhvQUPtVTcs5Bob9olYPw+hc7XlGSCZetiKzUMBOXXuD2hxW2P0BpyH66F6Ovuwb
1gkFuX7lJy8/8DI743VXo2nHJ74X3Pa5XcYr3iBCk1z0yg/DOndR3ORbwO8gHjLwT0beDITHl8x2
RJBNJAOjN8hkmI6vIZrmVlPVkC1zHCJyLrrwwknNCZZjuR4Cprc/D1gFWcqmscs3qvtHBbgSuBH4
4VmhW6cNbJr65qVHZ8Xyaf8gyR2YNsc2oynmJj4oRt/S+Bw+Dd7eRUfdiHIwlQqIHQ2cPuJXMEJc
DCDLyJSY+lVXFg9q82hLF6lQEiuEYkUE/5OCQBAkOFj+mPZk/J2NnKrGuxVVv1V/OWVFIfjFIniR
MfL5XuysfHGS8IdoyHr5RfldctkYUwB8C/YKCi/6qgq6PRhF8dVbraVFTdATbhVfgTJKCYATK86i
5km9cGVC+Sfv45fwZSz9J6JogKMbnw2sxe14EeHwnOWdhuOoYp+soFVnYnxB3UNTbQQ1mXmc4Bk+
/6qGVLTrn4uHBTUe+Nfv553gJlfMK0c+n2cwEymibiHvN0LYOlMXXjq3iUaql+/exnJJ86Hof3AH
LFRg0LdlMeBp8jsNBsaTfdWS0Bqg1g0fL3EKho222GHQdlPhBk8PxACPUKIPKDTw6RDKyoHLr7mc
qPRVi1yqssQRXHH+5NsM1hTkM4B+J3EbjJs5HG0DKGA3hmFgti9K+dhyrTI2AeFH2QLoi7H9yBFH
pbajvlRjavI9KXnWBnYkFDYpmEMJwcfPwcDY/gU8BIgexzN9zVrx3ku2QoFOM/tpJqxOduEcAgPD
RgfThar/UKRsogFsji8QokG1GoeVCX2pj2mGHf9u0nRXZRADmzrb6juO4bLtHy7nBb54074dgh8c
vJVH7EsKT4zO+xsGWNsNmI/Wqv9TYkV0380i+iHMXnlHXO1TyOV/9DiSZedFHjrZc4pJQDxalVT4
BKNyl5GkVUlWLpPJ70c9ZdajVloZIC+nGumykLSGVIXikr9JUucQUEwMPyBmuoeBcyOoEyMgNbK5
2m0DxDIGCkO+RIGbAUxfbGqvS3cZNmk6RNxvd0QS46JkPb/6csyUgMVocD0riiQiPc/JI9hL2scW
hzU4qBrA4eu4ulwlEU6GdyUx80UEACkZ6AF5/lgyk+OFb2KgAJKYTudBi2nZ8lql7N0o9zTfyl8H
cZihhqA3sHk+JLTWBlt29SFerpKkIEILNRp00nUB4vLH9zBFoyBX8hirLyj99lvqgBgm70FUTdL9
xyKkIRec2DZ51brcXf0u6cLiitVNbPxPtqBOB2XUcLXnTTgHNYHZ+Ig0RPbpuY+W8DIwC9O45kW/
VBSA9ECeh6IZxUyl6tQLOjOOZGafM6U4Fk3o/pthsILYTDiIVJ0OB8oDJLLQ1KdAd/A1jUbfgF/F
mCy1WNQQjGs2xYNutQ9Q6zydZtol3tnFa8vbl+2XEzFDx6ueh9aOmOf+c2P73b9eiZXSft7Qm7IT
2HbNfGSj7OgtfQKzAfO6+7jQgZd4XK3qwOIq/l44lrXwD2xx+EBFJhmYmjZNHf4lTuqdk4XLdzT2
/AtG3juvWBN7Huq2V2Q5WlytMADsUoZVy4W6C18zf6za1CTH3oSHf/jVs8ZtItjLCQM0dBFa4EuF
Ha5KabRDf7kO1g7bP34slP57NNv443vrl5FceD7GuQo74seIASEFOglxqnycNEmARjDTh8IfeCno
E1kHFbdiSV+sKL19aouxPHZynNQepLTsevzpS2I/axQz1eEVzR6cagOIKELGNMxi5bRiXCdVGZLI
ZRS8UzsEQ6pNdlU4Do7qHV2lhm70g+aN7VeB6Totc9BtbrbZqZFFmNuRPhOxVyAB7BrgM6CYRNou
9uR168nay0gG5wqcNRGey5BllKfNJiCq6uVWW1UWJK4bRyhyicF1sJQmWjyxRhX1SSZwLClzxXNF
JbouLL9ut5/zR+M5FXdkpTFSYdzWJCzpvIpRhBB5GdsCbCMkUxKHcxlJUP/0ruKC9zu2U7sK4DXY
D6W2Jf/tB+6znDnECtzmPuqaEUf4HyanegUasmE0+vHlUcRy91ElwBj8O2l63YjuiDoPtdmcgftv
BYkgX/gsStd3InVPKVLx/GFAr5+X4JTFmnNmDH5PJEAv68nsuv9rfhrSqnk+gLxxUKL3AYEwuaJh
V/xKr4fU8JqfxHARJ66xKhtdFOV5QbaMH6xRprcVa7nfacbO08cgWLxCD1QNdKTDKogb2VFweMe+
26sHk2egmfHyOgX8F/EzMolgjAfU/cBdiZTj/UEP3A1nkX7YH5CLKqTaGu/t/GVwSDUuy2iLUfft
ytC1hERGRo68oLao57LBGbTj6hhNCZNVr0hlF1G6xfUH70VhA/Kvjn/e3CNT4qN355hXyioJ4B05
5QUZwxoBz9Ox5rEoKqlzTzkkrx2h8ZxVYygDXDUHF4a67/tbUoDuTO7WTD5xkoXj2tUTpSX4IszR
9i3QyYFnmlW0fLxCbfASjBgWHKsu+cyRmd3IGp83U7DYaDUqWvAoSP10k9SouwCuxDL2jyZSK7V9
KsonlxABpzWTkW4SDNnjg5q32YUNX6cwe6QBPzbWZpOGttgOyA+dSBBgVffE+1oc3V2iXue5Eu8X
9ghu5TTocjIm4jbd995YfDHXxB7BTlqkJOdiooprtP/OslceWg6otCfo4wKqJKY5wHDKbGCko+uP
v6twpz7S0H1bPpe8Gny8JpBVXxyUFZxLm2XJ7Uc9IkQT1xMkM8iYYZSyHBOPcocowjgOIR117tS+
DT71KXU2JADeHS1W9m9TH0Hc7ucnMOIYbV877BkAOH0iq/FLy6sWuB53Vjt5wAujAfjtkXtKeTdC
2NWf6UepnKlWj7fWZwRXigmVUQHkgbb9aeC1M0LfVWQ5CiaS8yDntNdzoU94lXIXl41lCMBGlOxc
QU7jVcFXMIqClu+Bz6ateSDiqqfiqf0HJ4UoQQte68MD/C+1pD7ckoLh4wqa6SN8fzBTlhOF59LQ
HhjImpeYZ5mer0HqWL/opbnpO/YJ0gzXaa98Xj5bON51IDfmOSCZFkbaQoiNSP4XCVpcJuCTlcD8
0Tu1L2qGrniPGoptszfRrYS0ogB8M7GH7Aan2ofsPw4dxY6xdX8zgMC9FI6VksGWjcIEDRZn7sz8
S1k6QW7xbaTfxeF+tXmxsqwBy8fv3CBafxIFQAeRXyv81q/u8YRYOYL8RpK+dPJHuyL0/bhC3TWg
0jQLW5Lu7jD0GcWXjSAgqPVnIap79Qo5DYDXyWDw3I8TDeO0ahFKsoS+RkSIkvxkO/S8YeRUoIa3
vbswnXLn8F2+/cX0sHU14IO0xlphNdAu4MfN7YpMrK448mWbXeytScOFfBVWXvwxg/VE0oZs4psp
X7TqXYhv18cWHv4g012YhWREWuJZQbeSa3EKTHHkJSUI7kZ6lzZZz7HWR1u99tXM+D9HEde2F3g4
3mwo3Wqv7ROZERjJe+HfGr1h7EMLw7fAnW12NzCQ3yWqFdXje74hxAw9DricuIAj4su+fZtED61p
2itm+1hQhPw67Nql+2aVSVsJlKx+6cRhSGx8dqLX/YeM09vCwghPLgVL/SfOQzzsyGU53Vu5dxOC
vcFc3YfQ47e+Z96k4+oxWbmv9gOEBL76G1dGfa5GVsne/RZMCozsgTNeg1KB8bXaf+xCxWbfItKf
5ddMbdiKw9qIu77rlkvHF3a2RcsGR9p1dfgD5il1kkzRjgCBWBJY824TLLZiiJk685Mbgo4/zQmm
/sxS2J9WrJqQ+wj4ov+l5ku2Cz7f3vQCkYwO7cdmL+5eNKIyAXt/oGuRwP9B4IdsTGy5jg+ejMIo
m57K3uE9RjMgyNB8GmSpD5IAHkJFJnpiVGwx+hV3sjodFPbN/NOtfPBnF/xuHEsG2nYuqIlhixJ6
+J7lj8juIwxtOyN5kppnn7UAsjJs6ZJYtv2qm4YkclPRVp3Nl4gzXwZywF/l2GPwomd6F+KYdMdj
IKfax7b/BUIkqsIvJlSkaOF0Icvm54Vr58t/ldYC0ibrHINSdEyIEtqMv7OU3YN0RBwAMEm6N7Fi
3MVqikZVsI0SA9u/y6IUIUM5oKeYcPlcNYZTfcAMRLPDPW6BsDJc1h2IL9SHb0Uiu0gGGRcPW5Ku
5lbXHeehilmvEeQseNXaLM/Yv+v2azvG1yTyLrdunVBzzQdQbHRg0ldp+PWvGZn4EhyKf0F3+875
1dZKgDjy4I5z37rlHU1+IuIDFkqZJrI60IgkyRzMkrRUatYdi+HecZAD/lxhK2SNBNdLvWs3L9uf
AVsZ1wwelQ68bwKf1bdmC8kCXkHWvmKq7CNa0py9Vm7MMPmSTz3Pks0YjAet26lhopb6YNoinFso
W/LXRN2XPEAWF3ZaTaxJRN+i8xH5x5PQfKpP1LK1r56g93prLuADaFbaYjbT1ahcJya7VBSiO0xq
TYIcO5+dKszO9Ze8YjRCCNF9UVLi4pBBXVwM69dNF2nhSZZfXzjqD2s3yX9neTX3i5IfXSp9Uotz
oXiEc+TX2+ReGM1jIgVVPfJbrFnZEsUIdXiMJcelIWXxfBHkXwL3DO4wo+kN+WHdoqgalY+kKzhT
axAJEWYLHsR/SCbIhubAkPhwQ7tKox4Ai0SXUksd0D33x2j1/sFeYf5dXzBEyu8VmWxmNOXi+c8z
h3PSMW5SCcLSKP02EARyc45dBwsJwFZEXNcbrEcq7yQRhhBVWKiSaM8FiKsNNXBfnboHmgLJ7S0w
qTBgZDznu3BPiJaNdXSWj32jKic8JzzPwtcuSzdg7rULCfNeqm8iPffhumdAK2hgG0wiyfMgiv92
bf7nEd9CGks/qbZziyICqzx5Ei29q3ZwbL9mdnBw14I0Fur2SBbF1BEtAyC6KFPw5uVmsQ+/timy
yv0XG5alQ+fTojpRFEA9SKplDIsWQLD8g3fqYIvCjQhsmKcc7pvjEZWJzX6ud6nGyov9m/yEOuZp
HO1ow3qK8LX03JAoCwNpPJms39TsP65+2WUyZ0JvHJ6wQaR+h4eC6bBFE32RjCEjF2rMqFGU1SV6
pEetdupYy1snRxq4PwA+ZO1VZLRO3XBXZWlZU/lrInhUQFKBa2TOA04wXJiHO1513lgjMNf6aQR8
jcSIBWAIun/uzx7XRSBimmN5mjlXaZeTD1k8B8bX92ws7ccLCDpZXCQQBfUxV/DT6y5jCLu5HrVh
cTZU2vGERDZDnnTqO/QWx0mG7cxxkj6MQvkZT1mrv8gasiLiPrXYq12kOxbGlbrHczMamTCmUVLq
dozC+NLP4t6HcNcBtrPVyDFl6N1a7OfaRTQTV4lCpex2rr5wpFTnrh/vY77OFrsWTxmrZh7fcwkH
81yKgfryaNX7If6hEtOMq+Bnw7l1mgFhj0eHC1Gz+UeCVKqPq9mfoaXoM+czb1ee2HkSvjt8cCWd
lNy+ingaisCEJ9voXlKD1EXNlKyrB54cRa8mrMFK0hnIbwUYYV5HLcLDfNobzqzm+mZyqwW0ZANz
0HGjXZd3rKkG0bxcZg2AEZL4z1JFPDajh5QxYt8nOO7yXO6X4igWTSirOfAeH3Y6VNUSvssb0Rwv
rc0Ih0m9woUL7kqI8svhgd3insgADPcRmngLoOMpkC+pUeARxRCg8GewhtmoCoB72A6yGJD8zzTo
LKE9pQU8NCU7S+aq2BGXx2gQ5HPegtjr4un1Z83YXf/N7rHvD3fPFmRD9WI/g0nMEnc+SOSKAdhD
ERWq2YjhdnmzF5KEXdJJCfiA486M++RZVL5naK6tSBdxOizgz/cUNS8Vr7smXTAKRXZOSEHQV/Ik
wF9Vqp7Xk7SJoFzULmcr7Vp/PzIhL3RSIhitBeN2bOzCH4G+hZGR7pAfHLoig9SIq8ZfUDbUu0kT
vibV4S4H09+5DJ6zBdVZygvATwIutYd9HHTq76CUB1kaGkAKtCjEH8Gg0LVj2og8F2ji8v9ygxXl
YlhotnYSM58t+OBQUjB/rGaYEdmDjfSM09kTLtIC29NLS2fqu7XSGEhoCuS/bBKMo4UgvFTJr5ru
58iMQd/EMfya1gF5vXqFA7YxS3qAUw1Y4/zGLKABByR24OqYiIQz1kPcr+SMvotDFR9FLuJGQ5Hg
Ivr67N8MQMW/4TqZ5JtxXAkd2l20jSGYbN1i3yRqgTG1d+hEY/LVlN01ylRdv3ul30aRvQTv6Ecw
lgfuhVq3tbwQ02jdcPbflfpZpK5nbgxKztaerZt0omCXJKMlSjjaWLZajD/DW60SnIBBxWb2bNRV
U8fZRt6Ou8HjvgF1a9OL3jhvwj4CuEYGQ+fL6cTvI4RAwpjFJuwY4zOaaVHYObQ4aSSP3hCzuqOE
Xe0C8W4uuBOdNhRer41yG0/3nI0PwKeomASCaIHg4bkr3Qe9XnuzYN986nAKqjiODarg6oh8y0bt
tgTwpTxdn6TZ6IpOHmh+ECiWprD7tOEjzvGExmvu5cC+ltiFaC8Vda9v+FjRGNgJ74pt9bv5aAb5
6t77MCXg/XXDSG/LoZ0KvvsZ5UlqZQcZBCFdjATQgAZprmFf2MvO6EOxd0dtGTr93IzcZ49r9CEA
9+v8pQZwxH2Wr9sc8Ed4yhjCxfq+Ktk9Cvsafa4UoDdy6iVWVSWq6Rjqrn9NYuOfDQK7Wd7cnKr2
kBcY0+yzrYWRSfeUWjpApYdQdmXjHoRV/pcGiRONDePfyCEwUwRzWq/qESHfTsZt9VKNpWA8m56i
phAW3ivMjcvECuP7djyzvXrDs/ak8R0nPy6unQV+BcVA2omF+mn+wvgteXA/fp1wKm1KyqFak4rG
UTpd2fLEwd6ss3CYsrJkY2pzyLf0cRB0IdGskmjhkEK2iihkkWg1BBqXntq5dMUoanSh9Xr5Pjc6
WC5Xkrz6TqQp25ns2P9cSC16x/GSbGXpgjBRWHb0faUmr2eyPcPu3Qt22+zH4Tq7O2GaXh6I/K0D
9D1sDo2cuRzuB9nSDlJv3J+Kqe80/YGJkqjTBLv81JrhKwSTybjmXORj+L44ZZQYyiJJRDlF1zYA
r49TXQs18NKb6mGb2q8K+o/oOHiKsHk/wi2fGbO78toSQPrioQScoJ42Y3OYs1RysZfOTgJD6Gfx
fGmJaP7Qv2cknSrsGN7J5GsHPjJGGJtpunYfAiNtR4HDH5Ev9euIA8F68yGQ+S+NeeiGMdZgHfSq
UaITHH9Qsr6wE5YW9gVrwFD8gcksNgk3xoFQ8wtAxJBQGIBVACdU73hEIqrXSAj2OKmO75cYpHp6
87qmR14X3MKHS5yESmisR7x3qK13TMMbPQLdqc3Xx28YQ/PXd5oRaRlDejlCPFHVqlR0+HFPhQRo
1BpAgW8j4wrufm2za92G+S3Waf+6x097WomBf+f6hVK8sew0udFZyqQLxaMproLGFu7dRypqQcQm
GS1eLM4kIBV5DLxRhgBefyuvnK0EMwm1o2cdlKgHgZjh/xumg1RziFPcsgZcXWFpZIdQk8y3IlMx
XGKsWYlQn8PEb4o9JTYozjFiZJdjSLyW3GDUa9gU4//UrMwA02gsRqETgBHW9tfJ1tTxOYq7jnMh
PIKIj9Vu4+/VzLn6iEL0X3aywv/v/FiDLeUFVN4jzYjmt58/oXiuRN3/nIxaOvIJhH6+ask7b846
cWjfE18Rmr1pgt1bDVCOVzzpTJx7JklrERaI2jbL0rqUKV+rO0GQgCzPZ0/TpNrteqClYOgeKmJl
pXBoq4EccEuSUTOVnTXD2NZa/jXoWD+qMZvNPGUKtd53Qz+jijf7GAjtWyOtMcE4IIczawLTAw8j
2SxY/xSiYPK/LK/xAufwxqwbfIIHmc+L5QAr5Q3JnpMHstHv9haQicg/RpDhtiRCdrAhJhjNyzHk
t8hWLO3LXUnpSF5OJsPw5tpGXf1SmHB9V9JcpeetdU3JOWKkOlgotTWs0gtSATU/CCnxAoBQmhYK
sHo19DezLIdXWQyC0bWfrAkEKzg5GHwWKOgpgAm+lgVTToG29EiDOWrYsbgCpERxFQ2wilsQ5ymp
sKw0gxo81wjAo+QVN3cugl+VJV+7VZn6P0yRVxCAr9aRVPqRai69NXcoKJp5smaWD3gGBMH8eNiL
Vw9mtgrAQBL4ERfvrUiA8C0S27NaXznEDOl1/wGB+7VeRQjTr+GR7spbVFyufC8LS5xsYZtwqPZq
McZQu+7DRrB2yi2vuuCl5fJKtQZA4/4iovxi7hRfWCKcW/zR24AedKwLUVF8vi0tUt5Ad5fdma5X
oXgXEP/yWd9kYI0UJfyaTiVR/f9vrgqJzy3yTlDy+mGxmjHVrt2qKU3C3TEWUWjIFwECLeJpK1Wl
Q1zAcJJ5dYf8xTZiVHflvWOkktLQWnnJGw6ye+xJFMHrfUJY8RdDtJCVk4AgxCvnn6uEHTpSCncM
OjdyySiH6EvlIGRj1bN+FNUo4BqTQBonX5jxbI05FUJcPVhe519kvNMixKZlcsBOAtE0cEoMQ1tT
H+X84Rj22UQCheMfy/8JWGCUkWpMu+e+gK1IcefTAzvyCe/BvQGxd2RXqlKPnbZq4SsO2AEiqhTo
rFKkTGbrjE3AF+pLa3qSItqeZlGDEPjWirdnsu9hVqVFyeKSx6n4eIKQUi7r5rd9SvsnZgMBTC5n
yUgZdkA8CoucySadPFg5HSuPMeI2Q2KxsrlD4HGp3FoFakzvEWU/4ZYNkXlYQklRjiqdGOnxj/5k
QnmcMq8ZEz7M6H4VWolsYHFUvY8OYkCLhAU7tK66qo8GXM5nHf03DHNLoBmlC7naEiNDco/qYkS0
UuR9IyekLpnPFTOxbxFv5BH5tCIor5yUnPEhNuPeQAsv5AkqzgcvkSMcZbmBSgEKaJMjroYC/d34
WfKd46HxwPhKrJl2AI92w5PuKIyDZVoelIfelWU8EtA/Oek4MJWyXR8XTacChujFxZz/8PNqazUo
PSnpvxUB4UktvlBmzDf89fWVJH+OQUZBufcsbO8eBNgzFjvohyHjorldoE1mDm+Hkbu9CesxXjoG
8YiST/oVwqDeIhWtfulcQh2m28FcIJDmJDkmuHgEBIlu7iLcjizZSF2VnnGpxSNJmWIqSx2hmzpN
0yL7GWIP8SJcoJ1LVaA6qWIZIvJUp06FoHCvUMvZ3W8pDQrUfGZ1d68hYocfIce2jMPBtIxs9Xw4
NuBig+MY28h8JgWacLaMLqzX6lcItr2md12V7oD2fW1seu3tfyn2GrfLbHQWorYq19zRViGXxtAX
WZJJUGJyxMiJIV6UPqGBgudrTOHV5U6esOfjZt/Fe5w9EtzagrX7yhLpVN+kjxcFS4mYs2n+HnEE
8zm4Bz7MpRK+BQZWRlehhnpHIMMIdtjYdYZAN0TE4Q4mms25fLwH8n+l3vuaSjuwS/TIUcA/ZGCa
5/uCyzKErdmGW7vPMNJBJ6uW9en2M1Jzcrb0lXm5LZg/kVqR/mc2IhdYpFJ2lHzt8y9l7dFyCuw3
CYlK2qJGZC/bk+66az7pR+XY3ZGaAUtUEoX511fu9nVyndNbbVv77/m+ovDaLxRurNqctS62G1Pw
N7ZBP4sPB85EuL2gI163LxqllkNcXOliXBSMkz9Mxl4c2tW0/+pUmlIxQELdFmrhhow0R7SIAoZ/
aV5re+a7JZK/8j35QI5kZD6Iae0xGJg/SD2BCElm7FgMicE/SS42Le5WFCmxj9hihldJU5ZoGA78
rOhZZl1wBBNIBPRx9pmeZYtEdYINa/wOP8falzeXDd+kbo1isvPXMwxwZdQbYvjkhNlc7FhCI6ie
JQKPCaIsHjQLJmfXjZ9m+Nu6uhJmHK4EL0hnkgbao6UuVVBQlTnaYxOYjS+Gd1uAwly+QzGMC3jk
ZXVwa9VE6vqtUz3AnyACSFVBIQjX7jQD3yE34PXfEfwrw11bx/ksUEudNEe6LjbtgPkrp1gh45Ww
/45L289Cn1z3FgOAnq9cqkwdFRTkl6LxrdrsjpVIccvT2+8JUTmIGQgLLOLaJaWwwcSdENoN0B7w
wV0UjMemrkvhKctO2s1if2xhfaqD8KyYXYo8t3qRIRodAx706Sg4WpWZRv2FPCzhy+YV313QWjNa
OMsv3i6sSsGvByiN/ND2jnE8vrkdjKU/Et+bjY6uJs5MtVITCjs7hWNKhV+kzoaiSYNSQs8trGPy
3GwfOs5DiGeqeZhohV9YLaISEh2NqiDbrLZe3mevmCuPJ19Krb/dAzdENblsyhRjUlws5tor6/jj
JaXmVhxo6fEi5Wt/dfYjAQlz1EbT1vwjyK3XhdPiY4s71/PAUxejy6RBq0gv6EOhVR2YiiR+LLmP
P/41/e0rwmqUXdffUpYSHFwWZBNngP2HGmxWe4jRPRMyMmAwen1Wgm+4kOOpHBih53W2msP8uwd/
vSyYgCsT1Pa22Ik5NmK27SNZdpS0roe5C902LeGguc1W7moXXhN4nqu1+NxEy3r3lD6pXlMGyxJu
cBVhrFFM/WQ844s2qgE+mEiLIJOT0VTIz61+5ATjsrrDKXKCzkZhCtC5L6jPhjIdIMPMz3mIwd6t
dTp/U/lH2so8x4nCJ4gefPNOLd+OQaps19lNLxMqWYzh4nJLR+/TkMBPoyczY6QJVmma99x0PH21
IdlnFdbBLPprs7QzQ/Xld5t2jlf/QyQWeqERFKAAIh75WO23WBCH5BAmm+UvwJSm7OtRftODgKLx
40oQJMIlGEXSUcWE4/Mznau3Y/96psql9u/7UYWwoHGzcy1+lU/Jq9TuMmldHcFpKDCmse3jQAVE
OE2MEDNvYKypqwCwtkwMfEUOnS1dDQ/PNth9mGMEQE0YMb+MEFjs3KDK8PXgW99ZeAm/xew6T5GZ
TaGkglv1N+IaSs/UZOYxR91EFeJ3D1ihxdNA8TGt4n9axTHKhpa5GGvqmQQ1PVpwwYZnqu7qWoWs
xbP+57nhr+n8Bz6ZzwgHCnnmsFxWGBYP/729oFVKv/w0ogsVS/sicyCotcsJU6p5fwO7IfMNm8wJ
wxPjNp76QIgyI0jPxW1Ib3aS5DpGDJH82uvYuSqwN7t0x+Tckl0Lta8sAGMx0sQMqPBj/oGjD8sg
Afyoa0kGZ2czCc9nSXC6SAPFp1PWUfmMHAlhRC84KXLIA1bLU0EMNH0ZzeWkxT+OIu8eChlAo/Zd
g2V8vLp1Tu6wM1vsqwLg4TnJQccLGZudYhbpgp7ehykvYnfbYPgsywoKbP7Vqv40fCqd0DlU+5b+
fIWaI0W3sNQrwprwjBFScqUO77Uq34xWjHVvWmhq2+jieyXitNJgZhJfqbq7DBUaYRTty9qiBwzM
8LaH9T958wjumpSiqwjTwon/lglQBXMKNUcsj1MnU5rsrHrPpHmBW1y4jNyHkIMr5AV19ue4BJZg
BiH57mxyc0XwwZD91YEUDy3cS0CA96Fb9U83pRO6XabdeIh7ADJn7BGN15wsxSNSEx7wbvKhcTI+
aYOlZhmMaqHeJXHKaVD3S7skpnBhxH/gG8LyM3hCJ+48X7NC98QkUPMUXFSTIgDqMiTUd+G7X8DK
3tE9kV7iN7jhKZ0FVocrzsUbkUontR/2Ztd3aJL5RBkio34hT5jGSqISuAEJYi2UmEWF5550wjYW
gxB4Cv32bkPlKGhmVwkOp9JigW/I08aS6+Z+RngF4B51a1Gxw0jSgLk4gkXHL2bI7E3lFeGghL2R
EnODOTeCES4xUzcz0xkGswMmjw6RkjCaOg30Z6O4xGoTThiTjtZ73PgkV7Yqov1pLTw8yKS5L0Be
WkaQYqfMoDJ0zrb9TtotXEZBp/C4qoNas0dfUEQnjlVpdbp8GVTTrmB61IuxT2MgRAw+Vou5t+YC
pA90Qigwnv7jWCVuDp3FbAFQL9NGty+f0i02ALEtcOF/iT2LUgcYUTHMaQ4J8B0fTzWsxOYuto3D
JdqJ265nuqLC179etYd7pnHYhtPIY9T/q5cQdxOl7ebL30WwkNvC46lRkrvlr1MAg+qbM8l5uUdi
pCglEkangrYuoJevvhvywOG330Zi2LitHoBtsaZllwjy7jLq2cRhmOkoYSiembvzIFRzER+fjeYW
h/d+YAk56X/WTjICpqWdS4KzkpJHU7fGwR1w2zMuwKMM9SjAZcBxeldoz9f5/QTKMjk0iXSj5fpm
UClTdc3PqBmOXucaiQndKwUWQtJ/aUvOVRIo+nVPoERZAF9pojlJ22Pheuw7sdcFf76uPVKNl5+8
BDu28WfRgixez+9ndYxuVulnOMMhJtr+O0LzI6K9WrGItSymBzqF9IGznc+h2LJP70FjU3GZcDwO
ARxvoCDaQKAawuz271VFuSwXF9hn4wXwwxUxenN/F7H+IjFzJO7WIm6iULFZUJ0JErq5Hsy1hNo4
+KKyuO1QPpo8JGDnu2jbBB7ZkONZHDnDoQ6Z14eL7LlTJAQ3m7WiFLjdXcybGv/Lh2zEOlYy1+3N
bKk9ZrfjvwNEJsbxbermlGAC+2zAyQHAZuKR4vdhA5pn/9v/tBvsE6F7kAa1Pj8Qt1FASF/U7POz
fAh+9QoEHr4bGjFPnCWeEqSTqgIO+BIXDdE0MdvmKygqImgDfLmxdh0IuPVNAUL9FHrH5yQFHloS
mHi4Bo8cY8bBKUZtcbW5ElAdygfn2E9dVC0xC3ljC5fBQUeOxlCDrIdu5akkjhc1Mgj32789XEk1
gcR4VXl6QcTGqS0mK5NBglyxT5REkHcV7J0tW6k0qvZo9GjvyL076t11750FVosnXNx9tdvzU6wx
UbBG4iSfp5MCro57eg2HHZWXxl4Fxs65wJVWQgRd6ElIqwL7sZc8K+PuRKNfM6oBbFWDds/W27fZ
38/Cr5rEX34N5EFIf5wH3manOAxW5XquzEmCXzE5zl+DNkQXr2Vj2EU+SC6fAv8lT5xPM2Rk0PXt
gtDYIT+75vw/i5mUNoWmvwXzmbnYrG4OeUgwdwJxH0oVJQco3QRNTBqmb0BZChQ5eBC5F9KQm8CD
yOl7Ct1sYPiXHGqH5Iv22AY4KlAGJEtSpnIQpyN+9B105d/aHho8qKxkTOXPIVGjga4+z2OxGhP8
7ghxeE+KW8swxyvjcm3k53udvRiqmaMBE6uO6xk1mmNmd6U5T+aRc9E+PP8cr2op81iCXoNrowje
yfpsEtS5+sEyo/sRFPf9LG5S8zfIa3esyzWErrupybIoSP36dgtbedVj9jhBesY1DWOI+hEWV99W
4exkjYuQ4L2P7ldcOpnLYQY6i4j1TY/PgYCrI1orfyQivHj7Trl8wTNYKf4kaYX4xxsf/GzfzqUG
3swYnGEjCnKci0U/h8mM008QGD9TIkrr+Kowps9EPqb38Q1EQmLwTWs9KB6+obgC1Vo6O3YNX8P4
p92PyWIlmNyyS6nC4b6sugTWNbDKC1OQ4I7shPJg1On9jNxMharh2mLLeTBxaWwHpdZOY33Nqp4u
0iwez4XR5LN0pPiTq0zLmmnxzkGbqbsiX4Seo4nFjSuY1w7sC9cFldiDwn08PT5dVQSCEMa3rIeK
qNtcQ4Ut+Y7wpQnmo88AnRktuFDMASiHo/v2WclGSyQWGiyKYiE0QgRweUACNlcLl3Hb2ezE2ZVB
xTm4YKj7jEZcfBnM9RJRXTRCh5rggh1/0ag3kMGHZpuzjOzFyK4rkwOmo5WWOXMa/tT7xHGkWTRR
he+PLzlp33wNEk5zOtMRoAqTi4LWWov2VobWPx1kacB3K459IxRAqThOQXKbTVnMYm3xzngIFqbg
Xn0uUejv+RlTEN20def2aUsjC8XufpWKR6+Xu7A2HKvyrIvfwluIVHj0j+7HB2ADh5QQaRyKR+EV
BtvwRwxc9+p5Ww1+12jevBBm/9KkH4StW7jmWxK3z1d2TWTrXcBKqLgFtLDmwDHcD3zuctRLTfuT
cgakPzvF/6Yuetadq+1ctWgOL66BgPIsIFdRmtXpebdZIw820wig2E6hrgH4BIe41OG9Rnrnod/u
fG+avx07M0FcOtbBkZ4jU0JTAlWk+mH5tO76NMJD1zxSLXHhAyXZSCQGo4CLQzYymxm6LYNysQhq
gLagJl54k+Qe3hhe9SiOtYnGDd6Ws9zJXF6ZWw4dJxLGmBHAKpQblAv/+V2y4z7fDs1wHLHuxuCJ
jGyh6yhgbd73GKwhaOjYuQxAJgjN7qtjywLNLELqkUVR6/q+LGrjlVww/5VSO7p0tS7uma7IA7wg
DysSN44gpugYFgwbFDgqvMinkhuyIkkUOtaps41LiKmBTpm93QllVnEolLaRCHnooBEho/Jv7TPl
rn2nb2iSkti7Xe9kZTrGfkupc4c7pFX4eltBuZytFye4tUKI+de5FE/V6qvR+QndgTFkIzN+L70k
B8nn+yf6V5kNzWNg2NzEvJ2VWcSUSJkCMWH7d+4U9cEG5Ej2m1mGCeIIMawM9xMkEbCfszpFuhzB
5EC86x/7QO9zYNfi4D/LSMAYlZVa9Sxa6sbOzZn7BNdlOwXgrbh5Qk72wKnBHhjHe99SU4+88x7Z
X6vNQzmhTOQ8YChI3D2uBEYHjHAnwL22wYMGMcyPOXd+UxLvI0KBMPwhtP9ys2sMRwROkHsvYr/P
I4t1WrwzNXv9a9B78h3Nr92Uaebnm1vOZ/g+YAAIdI1c8WJgS74xnVxglTlyZOrmpe39Q341/3aO
lFPQtJq6xjjBjwvlYgQ+0aNTMcBKJR/f7uy/U0IC97ROaVrODbks1uvEWuxTiRGpz7wYxUAJrLR5
uZ+AF8ERBLNJUDw8+QbkjeJFrJscobee1IzQ6FeACoaaQNSCYdBcnJ1nUfkMHAepuRnIBmugbkXJ
l/B9GyiFmPHqs4GgXfsWdg0kBoedtOatJfUlqi1XxBIygMwKNeK/edHzakCi/IcYh5yb4wsKURka
m3u8qKhsI1feDGcB0RdvpMeRhJnknb/DuJl5KA/x9jJC7SzQ+xIXIngZYYpZji0bLMHsiGZuarYK
jDY2jA3hG+tW5xWZCs6hEU5wLUGl7PHPDPLjt1Hst4Gksdp8BVdiGKT85SZmcOuSgg7mx4tzHoCB
dqJSQ4aO3GP4Hln24POjd3h9Mihr9hdXheN8SPnHsIHzq8/bKn4Di2p6Hls6LMOrysqhPIgd7006
IuQh/AqPR8D4ftviqZCOb8qaTNz9gNfvDDc8p23IFjteIOmHOpGqJSbIzLfSPtECl9dFiPBo4Fug
b6cosWRhW9InrNY5ufPYYLnoLzlCLMsUBIhWmO0yYUYDAXDy9LiPB7j3+uLff0RWIwrxKjteEuT0
hvBvXRqh/7Yblw624xQOIyeLHIzmjT8NV87zKjyRALmf6hNjqi7JXyOU1VVzfQZQ/LeKgA2D1w79
+nTugIi7NnhsXO+3VP5w5FDhmpfRsXFTG2I7qCgbYvxWWkqrUVoIanSdzCP4JiV0fRtmQLONJvjz
xgA6dMJifFvzFLv068LjojJqubeHGdqGMHJeWHqImLY/LCDw6J73TujpJROBwc4npGeuuSALols8
Gk40gCkYovqtOboGFw1OgWQSn4F6i/xLWBPyHI7pnGIjQi4cbGCZbngBziDmOvjmad7kc1w35Byr
0yWg94k8hu3Dj875TfuNLJjBSV/Cdwu5xO6hVq8tYNYI1m9JjhSITtLQud8M2x6sGyVXBtPjkAl4
qeY6dZl4+W1ixEEIbG3Aw86jqnx67Jta/g21Ta2QrWKAsFYfw6NFjVAi1ilmZjIeGWhoLQ+5y3JB
hC9T6Fn4aJ3AeKqgZvliL1QRID/pKp1D+/ReKrjMbeY2tvi4MVI2/FjOlGI0JvKR2zp3zPpifb51
kfsqTgjYEY8tKeioMQDIIMzkctmGRD4s/xQobrLTvZDJ74DaTNZrxGQ6B/Mm7ok8XJ+eHsK0a1+j
JMO4r+z7qg3ZPqZWGRMiTe2WBookDpfeI5aoMdLT0B4FKqlbvOh1ylxs8l/yrSY59MkJKXt9U7V/
xIeJfhEZT6zUMAGlsN/Jf2JdJb3oS1c0eJaBWHQRxQuO8MWCYwDfeeb4bqzL8arv7LxMYXh+10Hj
owypwo+EFMjOGJQ50urMdTppfWpk9FRvSV0bWGW4u18BrQZEjWOQypnqQAzkayUvSpQeREO6GRqO
ln/6/TK3I4WzoZ/FU7dlJZZsUJephwzieNZj0AoejjjsRePlnfDECuF881mdp6V42zyuCsqEcJOT
Pmf4KMDcKRQJJeOgOgmxop6u0iYq60BfUSj6vZlJ0IONjIVElLDGT2zq/5q2jQZiUyx+e3i7GPXp
iXA6ySdAL76sMIlqQLTRMmaeiKfS9EBLGrEspYjCklbJZLeHlklPsXGKgM/DFZdHaYibRQ5UMY3j
O1b4PpJ6eTYKxw49TjVCc2aVO4XuE+vK2yRCLBgUL1Bw+lGKuqkPfpcitX886g6TCDjmnumvHIfv
+ajBedM/ft5WgZr+EJ/Vxf6FJUvIXVrLB0FhmHXXo53HAxEwGEGXQZLwUqomd3uoBpl9QWzupQ5V
4plnLotLQX1cZrPn7+Zv+VrgyasDVporBkSdLmlqxXt/E62sJ8EEtxUD7Kf+okkgBG91J83YTH1S
5EMV0QBJmvLtQMuPRvXfqELWdgNUolnuu2Qz+kuwwdfJRDaisn1rlVXjz5oxCYg9SfswsjzGWQLw
JUydZJSX9+KjN3rNi+Q+21F/pF24jTMiwRQosuRvRW3hm78q37QG/VR9vq0FfqmkwXFqdF/F0Gqh
qiTqhAYDDffCoXgSGwk2GPzNnpGZAj+KVDTQk8ttjD/pPaYJ8k39rcw9g1U6V+2joTb6K+jOcg+q
7nvQoVKQV/0Xn1301gqsltpeU38Nca826BHot9fR7/LezkKgSE2flrBzHArH4cILGQldxoVpkyVU
j623xxpiQ1nQQLCJLK0eUxb817vibnt98Fj2KSqKGb4jDiFo8X2lDrE/hVo664gphnuJDGdbSz51
8snKEn5/orv3pQWWi15J9RlDWMuGccyae6d3yZTAjoQIMa7dADPiZhUgcfJJ9SGiTzNCRLlZ2FjX
0lgv2a5Sb3Gp7i151CnqCZWuICj0RfMZXuo5BPl6uYkHs1BZSIq8TG2wVsERkgXdL6rRuIOIB/ke
b3T6fTmHqteCm64QTGd4Hy6S2P5uvZr++IuqQog1BoCs0n4DVpXSvCpE1epkTz5Q9wkSf9Ncdvcg
Yh0Smb/MIkp+GgVMSr8L1fgZXo/W+tDifro/jai/LriTdzzjsEBxCS1SGMrIZe+LEX/QyrpV9zTp
SYRyndKxisJRDAgktHO3WzDwF97dsItCGDS6m6v4/GtYkRuNCldTZ7cMH0Fo9vxm0diEkSkAjaId
pFL7GabM8hu8eKbteiIgJEPIhTix63JsPYDIGjuU89STnhoeCJMGF3LwR3vtiYfvaPQ2q1soqbyH
Q0vrHyjWf4q5Iuz64TRrDVLjSa5faul74MjDYei+HooyaM801KSONB1v3f1wZd8vuBR196LOlQjv
M4qr1xuw4FBY7cIZpzffU6O1EOlzy6Z71wER1+3bm30qeEn+m5Sm30smtCW1b7aQYDGFQYpZlC+b
Sj33YubDHvlNMp/MqnH4PMLhFvNRjJMlPkp5ESmvxKsPpu6czAqZmZMrKDWk2IVp4mqRm39rJuME
4aPK/w7mDUBJztA3W5MtOAq/dYvtx2370nBBwkKQszOq4k56TSjfoiiEfA/YUTh2ZOm7lvdfJ77i
YsW4h8SvbIkPLQhL7gQI5Y7IDJi3lhl+bQIMViC8B4XNs2fWhol/y/NYm0uF8OrOphjda1a3xKmC
ENssvZI/YfMVOOOvrs8HPx6DpHONojGrly0yFV7JUkcC/ytECHRHq1ZcVG2M3dH/5vfyfkMQu1PB
8VX6rFSUPJdbiga64nHh/f0Y9tZZngdSv13C6HWIv0TGzu2GcJ9uP4JdUyaU8D+GRAMYZ9vzTWfw
AA2nsKyvTLzUoNs5zaDGhDmxU77HJBDr9UtOoHpQ6RGE5gbTOAyUqpLQS65Di5OszeSq2qa3hic7
u9jsJSZUWG76R/jcenFVttk/1pijvYBmybEpvatrt6WoVK9p4iYrkA5oozuEiosjIzb53YE430fJ
I/FjPwl37FZ3pTa7aw4eQDZtuSjFXGVa/A4guhApMX+udGzKewtdoqELw3ZWkB5rfZLbuYpPUGmG
pgKW1UCOY3O7brYyiyp1Gxqemu5jy22Yq5C1AuXJSbCfpmItF5Glv90qyscAs8jhFM7brlJyOg0I
buUIZtJ6+EEEfmPT1su40dwAnKavvha7Sse9zgd621IA3Q1EXv0+jRhid1qTuhnWGx+BLNCEtNEt
4QrLMey6C1jTrCU1y/TR4SewUgN71tPxtU+ja2WDd8r/YCXJG8m5DY8HO0LN3jAftY7bRwU1y3Xu
ABCg3RCwCZSTrj61UcwWL5hATfzbfFWfhOl88qozTO1eURfCyt5aLbUQuPEUTxTdRffsm/zNodl/
iiA/zkIrALI3QVGepK70mC/hag5WrPmcmDelddIZ7sd6gR+nPYYlJr7cSmHGDzBWHueMUd35AEbT
mKQk2ksh7sTs+k3NhqBJrfQMSvgoqykmZTvIO2B0oeFysTvqewcZtOamaXC0muYTLhfNx0i+PJun
EWVaL8tGT50hDIvJIfswFXbHsKtu1MvaBk8JIr4Sakjy4NSprbP1P7J9a0JbV6dGkU69bic6lHJM
daZN4Nxdec2MNPR24P0wai0iGDIGq8uSGyZx3/k+ksh5otT/vyQkZCRGdtR7mnlRhjngD3dW9bDB
As5b33sIgslN8ZqmvR4NTEWqMOT8pPgrpmXxGS7Dt29ImMBtoeBRAWiJEDsnlas8TltamdHBCKGN
+NfRSP75WszRha33F+ClMnaRPc7tbhFhZkktrQq8LYovDEYwk5F4gXw870458KkCDg2jnn/ktk8v
K0Ex6qvJM0cMOOP0Ej+GL8RbEdN/FXgP1OZ/xTOIHXVBw9fmZhIz7810BMRSUNE5SiNUqle99PKa
Vat2KJssiqv1cOFLhRlMDNMApp4kndV2E72CoIN4fC9R6HP28ujJXg6n3qA4xvVZ3cAZCBxTBZaI
Wzmp+LOI3ml9Ny4Js08dNSctt1JBMXP+sDJJXgvBDz49Hnc/42YzhjOo8oCB0MsYYcb9xo/R55zv
xC5dAIR/7vQBc0lsDaeZuXBLE08qg1NyyAGKiUSAaYqECOe3eUDvTj6bMUV/IXYWnIeP/SAmvD/h
cxx9HgRsbi2ig/A5nxGY7JMDedlX7GmAIVokcBMXr4E6PhU4/CcxT16EJC5bhbSTCjGVCi2MxheM
z3Z2DlDSt5b5poThITSRPI2OGakPGabIY1KLWy7lRwKKVVgRE3sUsW3+0HK6kjxxc8si1lAA10Es
SHCE0bzS7xF+54tLGRuX9T3CCHkkKK2vF/lenwDCaEsnTu1AplcT5km+CIFjuBxtb9uEkbcba2aw
3I0Ad2UvfK1/jxwEApA8XXWBxXnIcRwt55c/Xum5KM62evZlK49WEX4XmtGP1SR6dtENBLEv7jBq
ktk68hFHpPlcRMcDctS/syJ8qYeTDUM+P+q6cXEfjahQXVGH/fMdD30apFf7HV7KdU6ipLHcE9T5
fRGI8VZz/YGGuFG35k4/MXqwV00BLEKhXYeCG994nf3JyhBO0WXA3NLGCg13uPSUXsI9Xqy+LMVj
SJK8EMc6gveOooUgxzw1sEspGzumsv4GKrxvynxgHnSscV68MKTvA2AtUANxSMFNI1DpmNpCHfkv
8A2chiWF0xu6UQ5n2Y3atQaKUjqPcOQV3qy3BWqgUJiFwwCz5rHbfUNoxWKF15vLc1Gb/IDQQ6VE
JxC/fJhzVI81ubQiArZlKjDIb/cwRekvCbN/pRvQDG6QKlQLHL+0lQdc9r1wafaR5k7zDbe3ZPOh
x+h/T42MkSNOn6q0m44VGeqyT6r0zdjoHkusuj8HQN95GwnWqE3XBpcKojklWFbOAK2bhvvrMdXi
o3nDBfAX4loXU6vjOEhUipiqOzW2oKbcEBxPJx20etTdmTww/F6R4kyP5Mki6E1rmCPdSNGciwqh
KYr08bShqRa8Ob0QFbAyDpxCEMDW/V4BkJGAaldmD90kS806Oneu6r8KVnrDNxUjWZnSyz3HGVPN
qR2BjibDBPi6uOq05ggef/Zm6VajRo+l3/+mvoR4WJyHMLNGnlWuT8WKy7kYCDDjfLrqhVmVRJoh
DTJHC2OpXgBttNqttfnsLIpQq/aQQPcN22hMlVHfN6qJxpU+gFzE2ngyPl5/vsUlvHCdW8mCnA/H
T90E+FY+Z/tN4dDG/n9NFO6Rq/qT0oV+ETO6sVLQ6cniL/XO+lX+eVFe54nm/yI5vwN35RKVbn8H
a08Kf+dv29ZdnvfGATaZSTTnBkUnj2em5oEEmj0feYNKF3l9yiG3e2gQIo3g9XZV7mg+y8iNWkch
JMjt6F2pcwZ1PIPrI1ofcX1BtYFalsQ7Hmq+KtrBmi+QcPUvu+7j+ZHk8okR7ahekurNW2imuvxp
pxrbWVrxgrDgHFwKUqRQ5kizhVpSVhHvsCis9+mu6fFjNT41ZSVvWNlDRpypTZgUeE/ZCPSryBFN
iDM7z4Xh9Rr5QsUhMQiE3e2FAjMfbM3Wn7IT1sLFCVrpQPjsujmajrhlUFUd+43rcAcDZfP47C+7
L/VA0jO0FQVJ1KOnL5p3SukLgjz19iizB6j12dN/M0IXLDU25DH5D/YLoENeg45O+dj8jivgT8pD
lxyYVWJYmiki9t2iPgZ/0CvBIa89P4bVP730NJWAq85otTTyH7yquJZ5r5v69iSeh1GdiMXY+8l3
gSpVOBZPer6tgkeqwy/wrHgbOWtgo3clqz4N4KmjOAkPBaWS6hdNjXmrxfHEfMHlJu1jvidWaQl+
28WLGo5+dcqxd/I30KrFj/jn6ns395lRKuVr4xJQ8h3GE2dQweYJj7g/h6NhBAkyF0pM0lF9xb91
Udyh3wUsRacstUR6D5lTtM8HB7L5w85OtirNo2NoDLTGagtDPRrXzQ8YnO/xgMhkwTdMmW0YGWlb
vM7PRVE5DFFoZVjuN0CLZWxGcRzKegTF6qyMXClm3uEXfcYkBiJIhP9zZz0O6vguzVC2xA65VaHg
isyHehK8xjZx7RKEOqIczpQ9BMWm24rAIFHoN37zD/9jFpw4DyPWqeUUJoTSKH0OtjgdLB7N7pf8
NRtuPPjB6MJDk4gGmCUMt2xi5QcHCSfNcgguu7xRSjzmB+q8Gmct5B6fHpNg2ZgFiRMmJQLJWS18
D7sSyglmWMYEaIz6LYc5AMBjZSoE0Ftk78OiIdnhLmcSJE25jxIAMs1u5z/fefWu8RJ6+FnFnKdT
YX5PSwGKa3LsxbqdJQYFQzX1GV5PJu3Ly2CsBsWOP6DYMXVn+BVOAxiKhkBqk70TATz9SVnEo1eT
gO27P6pnNPUktZDILSSPghk0ghzJKg4NqwL38dSzeOKDSNiHKxWQGwgbhhtJjdvq2JlRDjkudCcQ
tPe0cRzaJyHLn9QWDZZmVWVJJlkNLTqwXRBxSB8GhcLpQAt9xcDa4O6mo8tR9NLthLrwkcCJ5AUy
YZWzPojNBp2LP2JG8JMYznev8VrRrHPekPYDkWdH7ZKNCJC+iizbABh79v9AFgJSvQ43Bs+stuT7
mGBgpPlkdoO4k0l+XWUzSFfAnVpS4ykS/kJ36L0WVJAEeEGRo3AyB6L5//JCtfKlTjdhNzz43tds
OxJ5ymk2AKU99UN9d4hW2fZbiCOWC5RM+t4FUH2KctYUR5cOT870jNRkAeSH8Zb2EfvFQa60joje
1ZYYTj0vmUa+YgNn7C0LA1GQ2Mq3cPtZewRE188COTMXnBPF6kW14P3PAGdoL/g31dQ0eLJjjzRI
EW7XJEBOeaXUpVIwftg8DI2Dm5+iukeFSpTgkl8TrHgeJyXAFzRd2gMNoh330B6BhsdsAmrBGwha
OGJQwP5ToXZnqI/xbDI9FaZUNzvNu4AMXY9JSo0oZphYWDI6k9pbQcQ8L3sR7S2zMBjhs+DdqCnM
qKdxcmEeZjhOToZymI/ZkDVi2QZkCZEEwYZ7QObhZd9rOp7TsS/g/vxI/aqSinUIvQzPB6ub6atg
rFcJ6mATZIIJpLORh/ki/0WC/avmxTsvjzxNTwetgZ6OEQPerpJLe5It+Ya3ZiaZnB740TEJB0Y3
IHy7OWNl2ydWdiChLUD4krOE/xV10xDWw9eDhxh7P1PXenEOWnHnnyoE0bM2RV8Zer0Jeh/wBlTI
e509S27s3we72DgKcKrejCpPebIFL3I6aHy9NZlzLfkZFxwyFrRxM790hZ1zuYzCoMS0xjKsj/ub
4cx3KP241b5xK7lRJlwu0jWtCm5k0XYMUC4O21N1ypGmdVzk4gqP5q1ILOcbMxdyt0cLs088pX1K
hbIPlCJL2vtrJHDSTK3nfxHbsthNKw6/k74VD9292RfEWyJfac6ucBacgzI8XbbQ4EWC/6u/9GxU
0kl/jgV/acCrnEYgp0AcXay6OoUIIFZOkfG9ketQ/96whBynmPZkhb/mYibYA+Zfg97CX3DG+CX5
t4wf3b4RtiRAYNixoRrTVA31B+i+ptlFs+Jp9uJIO/l/9kkH8SDL32VcPUUMCXKBHs8+Ru7qVhTQ
vKjYhl1F9rdCEp9pMQid3ZBB1cy4ABoGaYNbZMD5MICvNtEgStzZpP9UIdWtdmZO0mRkItjeJbAL
a/+HnBD5ltFfaqEaDPS0/WfM0/BzMUOj+KaSL5QujhhQ7gD55BQAIwGnNvm3rVOHmjn7FIzz5LSH
XwjXtaOpMBUl9hsCcZ9hhcZEb3p+7D0csBQNBN9vuIMn/gH2aaq5uhn+98r1hmqH+xvdlosRJ1q+
EKGUCczkYzmDDrT/+fk5Z9tmRIzu5qeSpQkpw8KNlgPB8tHaqFrpQ9UTvmDCNB4U18TWMqJ+G692
x6ys0bm7Xkv8Ht3+5QQDZOChnsLs09veI2GcYnU14f5OiMezrax58pzMvz7dY8m1rVL0SPBesV6i
K4aVxJf4WgiAmlhn2p5/5ZB8PjVtjDG2mE3QgtzGlv6vtS/OlUzO3trifItajcrUsr7gHI/1lsng
HarWpbXcnngmtDK/JhcSAukga0MBoyvzav1hK/W8Ug2gkxQrc39YQe+/AWeLM+8tMMq8+rpu6B8z
WDG5zSQT3E28dF7b1f1Nu/kWpXs08crsfr7dvnol5VYnJxJ7MrE7C4oO7GtACKe3kM+sXWYdWsAR
QdSpAXzkaSoRNzImXMJL1BhcmS67S17OZ9ZTHJgiO3W2s1IuTOLnAdBNkQjgrONy7b9Ge8W36YBz
Vu6M+b64voX7C1Tbdx2raam/UXPH+i81iq/Myd9k6gHH/1pbhq1EkAqJybL0zlJtIwX7Kk6t2Xut
S35Vvi181gRJu02AIrX99++lw64PR63MV6o42U0ADPX7EWopuUXyfAonOGo1PT/8fcTcUJtLBymp
A84/cIoISD6pA9LeTHrtWfKtiNvK0DMmiV7+Dd1bs3csTNsawkSGKJTM83WoA46BDXnK7Nt1WlQ4
o37Eura7c6dOGQ6iRaJzw+Lx7q+hfRgWXq2dhFco1Q1RN14ZQBUiSdKu/8xM7LWVuwdx1pXFhgND
kKnTpZOsnwYU7hhDQXypt40dmKKbhyf1AiQ2zB7kKTIuazx/tMwrjrVPg3p7TFsi5BbJqkFhsQTz
hvrfFAd6cA2g+pUlOr78TtgYwFllI5FX2JpU4ZpTccQXuAOe3Rr+8+VispAIbl0Bem4AnyG01YLw
Yqq9jqMQTePGnH5eUy8Ea7rdMn35dQe59jI7/UlFlqLZqwW9n/o1w6zPXONhk+1s+wXJ2PvTS5lU
/zs2p6siUDIY4E6zg2BcsgVi0Creq6iaKHoYhpkBObWB4xjFG0SI92PM+TMpbBcJQXFpsXOjXm8s
Qs8WoF3MD6Q/GYKY+NzaKh8cdn0ytTb8sOPJWsGzRMlIuaakQYAtHf/sM6JbbZvRrw/HBc34RtUy
JxisilKegz98A3Fnof2JzDRLOK3x+9M7/Z7amO2Cate/jSY2hkd2j29rWwH/7pr0Eyc6cIc7aQvV
9fG6WuBJtSRE26XDBiCTdj2FcssjKxFjvAUB08BRWRGRyswhWw8ZcAY2lLvs0lxsN/iZDs7tJjwA
29LDOsz4NUhgtJ6VzuR5XmmC4pamHzIKkODxc6bIXovRVDxQcHMZqTJO3WAKkwGPNnKoGLZyIJhn
IkO/UbFLDpRVhxu0Xnp/R/R2G0sGgQIIr8FACTfAohZiO5A9k5+cncWv/QAX1ln35wtbU7rXeYYu
XNlS0I6XTIgMlqn411r1bViXmxI7c6COe3h+Z035Qc4Xm2n+6mrLC+CyiWd4UUDPfixz4eAykVF3
6zcZsBmh6QDMUfvNIqYPSzBe5bHcrCsy6LnpxKDefEyEQdZkzWI24AOxWhtMRhkjb+M24DKlFu2i
Xv5q887UBC8K9fZKe+8YzmkMCtgxMy49GCKAN0eKX4DUMrlLsQpcDPiHQILI6Dg/aqomVtefJaE6
HGA1f6Jke7kFfko5HqQEg7/PHuGBbscXwdROFBOAGBMnL5kpfiitpy0dn0NgOWoNNpCFe+NbCgfA
g7xYZg+43Y3RkLYg3yFl3Keo7PsZQMYpn0yBI0AgMpnmYt/zuoAADfYH+1yuvXvnhv8qf6A6OOhS
XTkSSvSajI7/azSalhsJB0LcBf+F7/kdZlI0kbUHWX8AZl3LxXysKoUH7eW0FGOJd//2yiO0JBbd
Qe7hfAX57hM209Rr3ZMrxBabxAc1YmkN52E047H0KYsEMsc3ry+RWc02gkzy0qaU366WmRYgYS+b
1XxP1+mn+NmF1uIJ+20TFpLfm5JsfozNmqIv+R8pjmX/x4i+wyp4EojLZifd3mxpoRbxydB0PKd/
qy2OQL0F4i/An/ubi2FrCGJVhyP0wTTCPj4toED3egEksPNtTunXV/J41MOdwnut270jL17ZTxIY
YzpW3zO248wlIiI1vzU0Yfz5+6bt09RdLvDvhxoAX+TmpJfwVdFVtmUAt8ayu5L29tK61OljuzM2
XW4fDFmmupdZxFw+LFhVTKozOfxd7JKYAqZyYLiIUw1dn/2cqMxjRuQpB1XJ2Ou/A9q9gvzkz3be
qqoEHq4+CzIwONwF1c7ue5ox7SyU+kNdbg5ELsb6kSNPASgGJ9vaO91cGUkqX2NAF0HEBI+zpzMm
B4QCTxEDxZHcEaYlGCIBrolZUJ/aoDX5yOBj4/Ew2nEWNsOCkc6vc8u6UF3yHxMdyq8zjT183xQG
LjoQKaHB232w3lX3rSfmSyP+0lqw8ZTIyEDz/9W9ybjyhsYtY+9efZmsWtC0q/dGD6G6OaFAd3hP
jZ0bnJr7bG8rcisEm5r+wHNET2ZyS/7pEId2u68mySoMx++EcUkaCc0zKn3sfUu7PY/G84YDdlm4
yKZhqEsqQHxHFICD4tdmtC6Es/zwpHVM253nrKLtVFkYLlV0X1MUEtkU2LGHfebJfXnLVvP6ZRNU
gajl5ekzqCo98upwaN6aGmz184DYBaZiCxwqhwkZZYlUnzGgHrWtHkkI9a24MbAXkpSyfOIUc82X
0f3P+QTR1zfzqsYK005EAUHjyEQPLSGgxylFycKeZos9VkQiIJiiXuEJV5t+6Wi59oA2euubGppt
gWg/k89fPEAkcpcJRDu5rnJHUVwVeGOeiaGi4hJ0R/6lzqk2vGI6EfvaEPehYl1QvlNC48sWY9Yy
146byhGq4/tlQpV5YaqSr1OCpHGsPblNLXX5vUaQd48i2Zux75UYu0tYB5G5bL+J/S0qZfakRMDG
f7+1xsrnTZFXD2ms2zOCIP3UlmcVESekywM/4BkOrEcqI4l4XRDCJ0pWy3ZY4qOrg1jT7e4rhH7x
Z4PtR+gMrlCDTWFPS07OEcrBzhSdehpa0yr4QXF0Y3V1wJTzNHMrUZRDtJQl55szMrkzUBu0fU3t
LIjlaDIok0ig7kSwcdPxs05iv5VGmRU1MdbweUEwrFWiw+FvInWud168R3bm7JabQs6dcWcneFva
pDSh8qZlAHvWFfsKJLk8cA1DX+EEgMg3CtA4x4BQuYJX8R6o4rO17JI7VpiP4ywYG6od6oRO0nJE
+9xmR77cGZ6k8CIOeN77W6ynboi6TQ9YgMXcf22F419B2F6Nwj3rHnWdXpkF/D0iHLPp5V84JQ2S
D6MCndZfSysBrItSTm3xwXNBnWxUR2fgQAnmCYIhsBvvsWuFdfXdKMVYwA/SF0B8UXztwGS9hpYv
iu1a2+VANE1LyPxWxjy5HytPeE0fA22uFKsHPjuatQn9d/Yr+c3PLkznQ7Hg+ExJ4Bgh69crs7FZ
qZF+9/MYxaEhtQLKT/HFGJU7TViGPw/xZWi04E6TNCQJiUN0mYVKJAxcYcq8udOtDxmlI6y4KENd
vM11laLluicjC0eKRKDYjmFUtpBHZcIX42Xq7q6BC3PMTiwnKBxsPs+TW883JpKWksmkLYE64Tpp
r+bGo1zF2pkgeOoQoLf0reyq9UgaLKM3hGj8CDBQCx/nvPg4LmjHtx0GAAxTtzmiFs61aX7BQozJ
vvApWd1fI+1nHxOr4R7KPqnrCk7Av34Yd9uUWHm4nhiLGbKKjjeKDqnUS61OIf+knVobFM66Kp3u
xeP2/bVd0CbmuBDkCFK7mgopyqnlY44DgAsNf0j8GcwsDoeSp27/rBvYQP/uCOpB9B+C4ogpxHqh
ZFgj+B85lFtCAHpe/Z6JsUfxHb3IMNcoRuxyxjIPc2ZRGZ4QZv/itBmS5xDy1U9M9TwvYFFrUUjU
1NFKZQVkuvJK3j8lE5f9r9zGXAWWHwgwKkQxVc34RhRsqsxcGCmPUbpeTnWNhVmtaQQXLYrPo12I
ZlNGH1s7OMvktftdxtDIsElqWD98hAomRZ0hS1iyAGPdtyj2nPknw48q//NTGNosvL+N2QO0UXEF
3752EHboIlCOsZGkIJ9kqMUMcVY5lXtwJHs9JpYcKboI4G+M450D2pVdQfjcLaepVOnDkOKd+Dfm
C1wXwSoeSSX0bNvlzVY3y7ntcxqE5Plm+5dRRbe8bIfVtOom3G40iW4xoUIcoiT9RYT/+9Hz/Xqc
zfW1sB0qIVSCtIr37NL70y/Utg0iE39o/MDbxRJZGmMoS7S7B1VezwJLW3roDandQkA8p4ZcH94a
PeKzOdwbL46fCQteDJrpKBtM7WvYRhWVq4kMfX9pZ2KKpffscUrolJ8Ahl6EnWr2cIrkVwVvCs31
KgegOjCXqxC14TwXZcEc9gWlCCwjCl3uczF93wI3jKy487Hk4QxalyqDsVJsVm0diKoha4gdqCjL
N8XC9EnvuyTp1BoKIx8BPuQzjF4x9SM6futPznlnF9ieLdMinSIip/eXMkOAqFOuO/l58/qVcR8n
kKSL8P1hxV56S7Xn/tnSeQvk2O0QH9c21Q/dRAOjbS8PLpt3PwCfYGQkEysX8bIGC/mNRHTDMEqM
ZNw20AlBJd+ISuMo2/R6qsvB/UGHRrT2JbNfKsalDn0F0IDsL0GVKaPqeEOnVLb7h5SQUzfOj2MH
ShMGVfTeIbA8MPABkeLb9Cu6ZRREldUQIBV0qp14Ssk66JQmyBExpCFSAphTAwBG6ZWgoRUZ6DTT
rNU1B3jBb1y+rMr75jqhDkrG4vlgo3pYlhYEC99oJCu+DXw+TLryy8ETcdLoxAycm4cAmXDVHMd6
cN6TQCrofiFcN+6xrwcu5aGsdt3QXuZC+UhDEqL7TeJxgG7++SOIT19K8MKxfLMxCIxT5EGHHaI6
4nYA5owaftGWrNbpqimnhY8ixGnjEm4atEEhNA3OyBcLGtNvMtZKQJOoK7j9u0GgGXTg5oUMu1sQ
wndn87OqLE70JE2uJ6qMoZdWt0py47hsWX0l475gXmZqJm5B5/dwSrCjPwSxJC/xq/w6H/EHG5gL
1kKbLVW6GYsqyA6bl/GMPyfH6McB2St2zIpjvyniJxkCZFhA86NhfDrQQSXa/1T3AbO1NnEE2xMN
7v63uwdftZaoE2lvuI1nqRBEh3vyB7PXAdJjXQOwjosfvbi8osR7ovhuBfhNISCWRmJmVGia5TSn
eF6ky1IW6DLMEDuGerKFiL+0dAHBX/5/nj2QDig3WGL6HmPzc7vaQ7Jla+CJHHxfppL+DmG7afuH
TztviuU4XErz1N/2fxv4OWETD3/+Oa20f9GDFVKeiimE/EipDEt/TGVHPDY0u1Vc2ZgWqxCl4k6f
fEtSXmZxe6kPDrP5QwfzVhnix3wOXtPPSC2fkBzKEJSZc6JNK8+3R+zoj3hslE2GxZCrDbNX6HD4
KkzCRa6Hyd2eCDUPIq4YZomZBky9aSskeQRAXk7dJjRV3es9TLFez5DBl8/D9TVIXDz3KhK4XgJr
oDJkZw6c24tBG+lW/vF2QKsY3Aoo8hx1Lfxttk2tqJwrDv8KoOzFs3z9Z7HNWoZA/oE/Zl9/eNdE
InKDIn12e7TsThRGNsjwLP0wu4x8++iUpE0l2iSaA4gYWW+wIQ3QgKJiyVe85o0Caan5RIRadbZa
aliisbPz3wB58yRKnZT9/Wem0DvqEExO+wGJVi2vylQXo2e8KowuSi9eLos2XC9gdlZWUZTPNqNR
3csY9gdcULnY25rrXvevM7HXBd/ubDl5uxWuzXTLlu48oSI5QvkDt2sJ7REBg2kGFiLsnldNQkq+
v3kwf4BWU5MZ/oCbGe5joGFrTF19ApoMeH4lq3unwLFCiy8ofmCmaxB97cXT6nAKVPky/GWVWFFu
SS5aOpFpyapmv7P4KXf5BjaypS03jAzzr+21YBY4NEnh35XuK3MgDurHvsl+odF98QW51T99Tard
DdXdItGZdxz7Ck3tBAvLFqH3Kvj9lfFVYMKRmPKZFAQvHfcysWYIaQoiWekmbq7+5p/m9R3PcfRK
KC0CDA74h3twYKVxTTmOQCWMhPIQBAtNkNBpaPuBDsd0MEVw6N6626eAPMZ3VPzyHCQm00nTlIlc
crvKXeA1lG07/B79lv9yw3FuDAoNIiye4GzTOUSNm5IBXcHNbqd8DPK8wuPYnu5NbX57Pw46kPzB
r1HwD0PVz3ZCU2PuDrZkMHx6jhzR965JpXJ0w65OkkKx852iin2Szh/oCKuPZUZIreUYdWmQ2kR+
7JdvAsg5IV+gzC21DO3QBtq1q5mi8oQNf1xgKHKw6s7ESw64q/YNJaDlcCYTyGTEgTfkAliwyPds
4mCfWFNhNGeqA8U19+OTs6Sm5b3+QdAB0Uvi10q1BH/pujjZczBly5iesOaSXAeX7aVMcvrYOZZR
ti9ws79F4VJodWdGuyTLneyVS9jNTMj5Kw5zsBlM+1Va7jxAFmf2NvuF/TvaztDawFFeGlMVR01o
Vxx1ylpC2ggwTiq5KusyTZ+x556v873WcA9GEWP7nxv/BciHY8YmIlIhzbBvSk1TgKPj7FRq9gqR
z8AFeFNtnhzqMO51TnK8vqsZmCTaGMF6JbwfbMijtXLEIRsPKl3OVyqi25RG2h/MlU4EbDfcppaD
AafuqC7AMsewIeIx1l7BR3ez9u2THeIyg3y8x2knv7uFjHHxY4GuUurk3gZMvguMnu6BQT6JBnOm
JywHDbZAhynBHiYftEYIP2MwmQ3tjDGhkMEStNYOvb7zpyCq+hAMjY+dfQrVyeuXMQXTyq7CkPyR
LKf7+zfAQeRqraa0Cy0yF0mvFjpuNWIa6S9XBaukHtnY8SwlQByo8qjetJcs4E6O2LVOjue6dnxx
NB2g3pmhEy0pMGMehzytz/xhaX0xLzxTE17KR3SZTHYlqZoPSPcPIg8JkiGslcGVud3s9A5N8opk
TYZtgpwe1twx0Iux5MmJXDhMiD10jBCq+VeABgJLyRQ1cAQF9KFSd2uKHN53tMnMdOMFfN89vpX0
8WsTYDS9irakgkHWIYDn4yFanK1PKQx0tGT/AJgfiKUkab8+UDGGboHbkCwKY6jDftjRy7OYYYWB
vJQ023taWNdvpcHLaXV1g5frktw0XAbjC9U76cHkmSQcLWsxMbdS/PaxsbekuTar0DgYHm6pvVND
nE9OWWvqYIPMBcHDaIpNSJAykGxop5Of8O9w5pIqE+TR7+3adgvFMrw3H2t2Sb8PCQai+kaz2RCz
tjo8p4VoMIbiqFWJxBGskDRZKkIVzPaloOwMv3sJBr4KwZ/eMem7r4smsyV7Gv/qveHNVoJ0aCxo
2QtKzDKRCQjFQpO42xe5AcE8OYsfTGloZOcPCaFnqoLbNlLr+JYoTC7EJ3TvnEN6QpqaybtazOxh
w4iplm+Mc3I+AGUvVP7Uk3+JZY7ywsvzgY82wOinQUwIahKZNMqUuBBYffk+RAiS5IRmpqRg1Kt2
tq3i0ZyzBm3MfLfmqTgPFp/yO2swFsA/rOGkEdwk9ka6i/kF8NzVme5jS8fodsB28GCkhnxyGm99
qiu7TFKl10nzQr7Xejoig3El1biqY10ubJ6gxoDY8063Koa3atMdyH3nExUsMTYcQK5hwaMmO7+z
eADYJlDBLyYbOZxwVMcdxed7bVFBqDD5JPfBOxVV99fEjo8BNOyv1cj+8iJDPPmxUDwccIMznMh0
tVf+ujuJZj22b7pz7OESqSb5QFRSy0XfKyVxPTfYDaj1x6N7mCGruDUcS7C29uo/c0BnPC+Of0TP
lW+pqesYCThUN7d7vP5w56eoHkNntvhqcjap0BI6XHqc0OxIuR8hLDpLxa4kARxVNNCMTpE3pHJP
X245YESKcnME+a09aIRdrA3usNVEmmsXYkH6fMivU0iwpSyk/I9Xv0PSK2HJDBO2qRi6vpUXvD+6
X1nBCZpuZAlNkIrin6/tV+GhLXC7mmBDMWqWRlHclpWIZp/O15QNxvGX+Nsecf0CzDOq84HXV1EE
E1eDeRx1JULdcjHvLH14bVQEp4poVh58YmxBWuWXfKvZpQEgqmD+jUjSG0tCrNpJVyZMGXFHn6Ot
A4/J3cwB8qbtBFi9cIWtbjGx9FqukJWbM4l+ZKNlCMXbQQXl5USdtr8BohM0xlKn8Hf/hyXVSHUG
wQ7pwRPmCH0ThAFd+1ppK+vv49LEP5Rpi85ZLUkJRdE8+eFtdHcazWG/Jq19q825miez/J693Q+I
d07q0v0QXdoeaEcl/ejcKc+QZ+/77O+WtHjmd8/7PgWrNUWcLYAdA3m60yv500NSc/fM46frG7mk
7I5ZYdL5wrpRvG0NJI6VfJdxcmxJGC6/TV09W14D2D0dX+o0NNtRbthMD98rtPW5QQhTNZAZ7FKq
EEVqucSaPF81TlrW8SbBSk/9hQwRrwfklUxK0COku64B9wDUEbtdIpTVdWmpOT9WabY3Ayem53FA
vE6PPZqQYiMd0k8JV7CZTlXzhFmTKk8s//3CQkrm8L/F0tmrtWFQ5F8xH2/5bHEBMKOSGGMvFd3r
58o9QOOvN4i2afyKdr/2/k61gTTmaf0EDo4AkzU9oNKemjIcd4Y7Fr8XRrtf6DO7W+mPB5TBUKy8
kT95pWDLv3cWKmpMM36aJOKoULJUZkM26dk4V7mwDJbb3NWoSnt1PQfZJuyQLA5MvZCOCFxcDf63
j91zL4ThG2HtJNjdUYvehuBk0i9IJHH5N6YOANNUp8e251Jr5BloOtThRivKOfZlWYo1eLu6xHzE
cuAX4vJ6mztK+bq2Ga8Q1wbffzSvWY4BRF3fDGRkvFg45g4WWE622wrbP+PiroOqLzquq0s0W9Xy
xsVdtDptAc82euL0xsf2jT8JK59O9+lBJtuw4WByrr/0hmyPgJOHFu20NFqCFsadFoidcr9F/8cv
fr4JEyN3RPAi3vIw+u6xsgc+do1xbLFzJ9+TNbg6Mclx7qmPOeDPJuktJ+BtfK303IPoiRwEeRxx
56ZNIrxE6E57He9Dp0THcc+eM5K9UTJfp+DR1x7VyFi2znYO7xNHicBe2PdnfEkKYoRU5gR2Vjsj
uExHd1Yn6dn8BXZM+p9kRGfEEZHS4caDBv2RDC/eWt4dzJriJkegh6qP0OcSgtIqFkGvM+RrAXZw
RGvWHGP9dStugy/koCOA2HZCQ58iWcSL3Aq6Ys+CSvGVRpcSdZ6OoFSmbkJGJfINCczecuq5UViq
9Hjrzro8G7dnfFawQTSSoIAQJFPmxvwD8G1/bLHYEZHwf3VXJfqV9KNZz9Aaqn/YJuvP28mGO5VR
vaDK7qsGSuOUTCc+en/11dfdyiBJeNlxH8YZtfQ+jltRDhCKwXVjHwSKwvmeof5uhR7jzEjIzf4F
CrxnGUkCmeGjVAH6MoR4jqRqK/h3565layMken73looKs94zuaO8C58Sw5CIeU6xWhscyQLtCx1E
Jn1ZlHEwrdpIxfR74P+9lKpu4FNX/p44QcocV4CU03qHQn42FWqcH40KHiZEKc2g5WWefnIqOTh9
HH3XNqEt2rvNH9/yMqzseLanJKUkU5NXG4bvngmPom2gHYBg6ycJOSC8W8UmAyuuUmO61FMcPAba
QCxeOX0pEk+UQFW7p2BPT5ErChFkIuxNyPDiZ+AtRT1QyzifpqlSQJtSqT+uYpuKpsh2Y5Qu4Q8M
oZ5UcwWRlkxfWz2LzcX2w/D1s1zp6Py/T3Xt1WVPeNIzKc0WkqJab7GPc5tofLDLUl985vxX0O62
wqc8KSy2wiwdH9wzMa0EjfKkeSCsD4hSvHVHAlw7AK86b3ht8+6of/IJPlDHfo5NNmr6ijeUiJ67
JAI51Bh72M+Ls4lHmCyk5F0mBL4SYZlmGCW3T9QZeS1sEjVy9C+dNDyxLIAjfFvoYOIDQmVzZv8k
AIn0NZfGBiGbTHDwS4NUx501KDkFePgIZhI/Nk9Yire0zGTIdqcxG2sBwIYvjh7XiM51toiNF/2x
gJzcDpROLYah9PVp5FquPeNY+F3gIf/K7rTVX52NoOXr89BWBsF/naDkL9r7RZonLqdFD79ppfPC
fQMl/ty+j0u1WTF/OvLbKt/lUOmzJPfLx4w76KXamjY78t2pa9qWCMroqy1/IQ3OAq+9T9Gr9D61
geM6voow7FVWFx9X+6Md2YILaH8w236UW7BGI70eFbEmHeSJny+j+V2cS/bbxDOhpsmp947xWPb9
cWWe1Aa4e7eXqGvo/vaTTMDtdwu9VdRrd+42OiHN0GhAsFcXBCuY4PYn9tTBB4YmkbbVN4xdXY7X
GSUw0DQHunK7l9q5uMtM0CfF0XOr82hGWxdBYggjz2wkCPsr+zv3rBXBw9UY9XISl26Xc0a5UWpO
xW2ZqIfpR6RG1k07Uq6KIUdx9tt7w9P+6vahi+F1Lgkv9gnnscwprdClmQzJ87FpWSZMcFVXkhGt
y3FWw0XVrAevDGe9X4S7V01gh7yV89YOdtnhJOX9Q833hTulHghS4QPX3XKUl3NBzLoMAggQYV71
WjdNIbFjcYdyDMXTUeegCqhem1YA4NXFAlpFFbzBJV3TYTMzlBE0nxeE+59AX+ESoum3iDES4bce
n7tgKXA5WJyBZCrp5t9Z+PddqgqXzZVanrdTYPFErJgZlcdA62zIGxNpqCi5R0qb2pB86KPpHUrC
jyMYZn6jCNjRDke7NrtqF0NWkoU+dND6fhCKxtgdZwQeQwGAnDpksUj0GHzG30f8XdtfMrECsnJN
Z70u/Qj7LUl+PQrKzZEm2Tz9NV2rKUXAb5RNC5olnxGjfhkur9YNyyjpcp/McAUbHMtg3tvZF8o3
M281ir5+mPTOOiNq4DusRAduYjIyDc2FHuDRLFbfbDPsiNHKcJ/SaVAbid06Y55fUI5Kolbt/x09
x8SxZh84pR1Ymz1xeyEqHS5k7nXRftIEo2k8WdY9a55Nv/+gt8aFpHfr6G0J+lwCzn7Bwr/IWICz
XUJ/HEHw5U6S9MHJPDC6aLqr1JUcEF0BRoM2Haj8NvPCPUIO3/jHibNHbBewlFU1HyEvWQB8fmNo
9kDUpDUI2DlLNHHH9ZFQS0imEfZK6FG+JAzepYYmcRdhuP1zaGP93mhNZ0GnxuIgrX4cgyqoSJ4A
2JuV59WtZ/7iSqTcIe7r5RdpJtr1QR57rijnvEmoILSfa6sk/DmG82zx55YT9LJGtfyBzfy4EBvc
0ojcPCdnTt1aGDw2QGc7eldpE+D/ejJ/YAfFWS9tU4GE9SUyfPohGcRbijopYuZXh9MwaM306tvO
IElMtP0+Gk3cM4E7jPLmnvxB7abRYoAxsEFBgWKdAT+1LafFixrra92t64fhGyUBxj9K8T09isId
E13tbnRlINEHEtbkCcMFvxsZ0zVGgvMvAYDeAQqV2tB4AWAh9bBXQy9186Ta9nLPxKVtziLaeDQJ
+NpA2m2z6HLhaa1cU405/olbH1T/OHLYUTdjhBu1YAgmPxeMzLyJBcg+f6YHLbE+Qg4WaX3ZXpT+
3Kyuh93NFDfFk6N3DfijfQwm/SsubL6tBux7dWBovmcKND3zV96Jb9uZlnUEA+M4UbId/7Z6IG8+
O1VdGlPoopWPWablo0wR9mCweqSq9UUHgNoICXG6FKLR0ZdqXPNtBYpXNkcrHWhBVigHpodOZKrd
u6zoKP+81iiK81/bFfwcw/3ze+PiFx5EfrXfKIM/ybdcxNzlYV/TlrTHHoN23Hc218TzSssRc4yU
ppMN9Q3P7lnnYDAU+VKuksPCKRDBmW22i/viyXVXQIfL7EE56LwpGpu2iUatkN1mU5UwYHZkEUxZ
XXHj3NRWLD2ZXRGrdiYLxZmA69fYNmOIBKbNv79gpQSSbvF5Dg8mGqrt0euX2xlNE1zSp42LQAzG
GWvULXf+/mnrogSrtfrF5BDeFNX0olJNjxc6d5mk9fp+OjSWjN8+RrIotk0nBHVL8vaRjsslOz8a
QhJaZnRKyCP0qppi4Joum6b2DaiKubpp1JGG8w5XwjML5KQvr+IbPZa3Xj3N7gug+bUTCETiyV2c
K7cHF8E2i0dsZQdqeb+bSF2tyGjc6clcT/6uBnDegtPFImO9m+HZY8ZEnmQYG95KSAY9XXWyC0j4
3LjaiZbs3FBIMLDgwk6Br2Jjg9CGFg78fS4UYusGrMlJcVy4JRnR26bj47sJooc0BNqcge3orpfV
qP+GoUAYBzPyk0O26zuyI5PohTgHq1MtbA5JVol23ujF4GGGebiesspWU6PAmRyWFtr2yusIUeir
ZghrWBhD9olnqZ6R95uEykKs8gRdR2z2lL910GqzWcpWcHe9OCFM2vmJioNQJ7TgPOcemwsF0cnw
kAyNVFN0FPZ10MJB3zsi4nDcn/Z1Y94DkgrJ40JAeizIDCffAITDA7wl66HO4y8eH9c8rJ7Cf7Sg
0hho4Y8RQ25/+EHTCFh859Bk2BwFJxF4orf3JNSkRqyH7+KgkBr99sf0GH0oNXajJXcTrQBCAuQ7
d3lUMJEyoJrgpWLmXyXBvDFo0S664HmXWFe7Iz14cO+Rx2xFop0DqDSeIddpQFVPqGbTHkwRUapG
D70NpKfySVrCm5arCd+hCpQD7i3GGd0tuf/sTE/VLKslMCR+CJwy35WwRNwNSMYkLcFXjAsNlniO
inN9zfqj2BUzp9fKTOQ+ovqX0Nxawze952XYUVFwKyQ3+eOJCZe0Gy5rEVK4J2LbhE+mOM+SvjvJ
zB3VjgJDRr1E+dhwrLvjRtIBI8+KtPpd4bsoOrKDqhiZpFs1JOU0vmoUS0sUGUjwJyc4t59M+F3s
C0nKp92RQ5yZuNOtxaZziiL2J/WqCN54cFAyBtuQ2gqYTOUA/B3ASbFKww7abvt5XF+arbPlwEUz
rxdI5Y6PM4uee903J6cKwdpqKvS5L84qRfX2bnT0MxQOZYF4omPpweFxP1XD8HyDIvABpFSfJF0e
E3ARw863tai7++jmeYWbI96GyTSDfJxHy9rVkIcZ+3eN8yrfMnUPVeWcGrKBh2xE4n2xwNdQ/x4n
EqMLSUyvvr6k9QXRyZh937ezNq4YxIPVRWvumBolmVWlY1SW0TvcKwPxwxNH+BQQExTK2WTL74bh
mwvxro9l897yv+3sQ/Im91NBUmOdksUFYeZ/IsCYjH8p20b4K7LP6h3pqjCgIwVmfRtPqQKXX12A
KleUjr+QGyz+8wO4GNbZb40WpRbmr+hVlK1w1DSm7qWhNsJAPP6EAUZgP6Ny7pbQQzkn2+49Kjwr
zK9c7LLWR8+9ERfwVhGfpErrFSebL33DNoMb38p0c6klyZlW9yOHr8dGpKNDN5qwnfBl78/kLKsq
kMzWc+mSMb7WBwYcxnbx7SZxLRdyheeQg9X+mDaYTg76lqmeKkLh6rTRMuaQ1a6Wax/Hi1a0E29/
HBwlo3z+FutOufYKViT4II+0EOi3S4zR+EPh5DyMV3FP4GRNzZ/OUPb4m1yBvUpn13Suo1z4PZFd
jHz8dort3dLwCn1XllNGpWLNIBL5SpQ1YLuOmWwapHfXUL0MaBsUTgSs1KcpdCocCIVSXU4ugV4t
7ly1Yyy0jZF9dK4CK4AosNGqWzvp6k1dE8Xh+r8UUNAB//+8vH9cuTEGMlAanIZSmUoG177ueo/v
0Kp7U9DZW6NNZZ9u2G0SWfBWJtkzDtJWpHPDoNeU2MyCCHbn0K/p+emJLHDenKaBviJl5/7AVPhs
c7F1X5BodMCSV/a77M9wLpvLG5fwHRJoEPZgDxbbk/sd79wROHMfWoaGsV0jKFZ3D59/rKnDk24q
Olum/v6hpGKpym0ot1On/MNLXxakqlg7555Qd4d7JQgb58JkTLj/RCgPVjsYB2PhqfvPGZ83DQco
3plQF1bidks98h5x0dRimLwt9C7EtqlowLPLK/lKJSrf/8gcxH6KtL1JZIYdzHzT4+j/hHH23Lrv
58Z/M8GgEoe5bJb0XbX4l1kd5QPsfpdMDGCl6/5QG6eMhwJPT1NOPrPj53gmJKEG2FNcMs6WAEO3
BcNCHLrNKHUtm/Su/8v5+pFm/ZVfSO+AIJnuxLk0ePyqmoA2PKDSOJ3uQKqWN3C/Ml5g4fINYs14
6jOdcKzSP96eXjnuQVQKpcQbY9VUnKWon6IilKZ9/7kYBl3mh7xBwVru/fha8v11Yl0PaI4X6Mgy
dfxCbrR9zH9ekhCWnQp6UTSHGD3l9J7pUrNA/F3rbZtAhhSY7bJCko9rBGId6w1NaFou7Y8mkXCF
dUzGnzdwaXoPwlsXV3bKlmhYuK7PHIMz5nnsp7+1C7a3hlFgewqZ4A3Epuz8ITBC0oFeKlrxWLi+
TGug3dGpkv0c8Ize58DnPLjlkUiQh4UD045sLmdjEUxX6QrEphXF64Z2okOXP85CwD8swVa5wKCj
fmpHCi1Vbg0cZfLg/gEaQggSpYSUZEUANWLZ0NFN9xxitkSCCVgecvpQXMCjmf/ZXRc9MDv7l1Dm
LcBHQT0S6IfYB3SZ04j5b8KTN5AOH0NJahZla5ZZPLfcbE5u8QHayWX8MrkQNkgcwMaRk9og7DQi
5udl8vXEgVKEOguPKXW0/NUQc11HQBDkqsqc5NF96rLIN1uf9WKRrvIkDx98b4PfEStb2QvQTDCu
i0jMhlA2sz0+UW/StgWIZnb5cRUcukRA4o764B2DWelxWrJzTBagJFSJFzVnI79vQl0p6XXDLHJq
KSYWu+J1EnZW1t6PNq08S2cZViZXWy2gLHPBP5p28NzrdDMXT8VX7mtui5SnxtgLrGmfJA+YWVUy
NWD0H71eCu1hw1Ey+btVFSaggD1VOvZL1/ojJymM4o1SvwGKMNM/jlJ1C8iiBAfGEIBSFHP9E1Tw
Xm8j8+Ke2jcS5NVc75kt3Q6wcOI5hLesLS/FQwteYOpW9S5lDIWHZEH36SursmHsMf4wz4MeGKKL
vjwp5H79PzEHFn2F2+RJ7sqqx/t7ncwUZ10QGxF+HmAKNk1ewjMMT2JEV21gKaEEP2t0Keae1Oug
M+f4YJ48x9zRWpzhbZgp6oW+2O0fVwPs5EK+bSTXcbvDApwP6SsImHhvWtSggpC7S563y5JS9pQX
1e+5G+ZYA6qPYCymfNtigMRwC+xztJC0VyliRxJy4Ffmx26C4jq6a7iS7NHHAyQFW0P4jKFs66eO
Od6FbnJ9mKgGAdzbAdhHgJmGHZM9vdrzmr6TVb01M6o+hvcB3KRMHVG7KfoUxPqh5svZ16qJUFKY
du0mQU29gLwZvBjLISfC008+40Zj1lXch4NDQHrOiMb91Bun+LFQMODlC6salwZUYPyk2QGcEYsE
f/Y9j4/tj2igWnvO8t4AYnXeRYpD0fjfLeiUHcBv7CS4vugpivVfKT+l88/WXIYF71n21KzOnSIM
a8qDiQUpwXRFdsu7dRyKqVLCKAmD5NqtYAjBIVZHpEm4CTvaBd50VB5q7Y3OZ41nZKHRGtowKn1v
nr1RdnHqmBwu72ZG+RJQL8S3LQTW+IatSMSLJysJ/N+M64vxuepIycTRAmrkjxGfZ/kN7Jaypu01
E4DaE67Ss3A4WDZu1WJAbSpAfJzjAYalFyGZaZMj17VKrdLnGkFjqslv+7BmdA0LbNo43LYq58ew
QBgGMR+hgGOp9/HBCWRM0JXCR+x7q1Rx7DLZm7s1sXJReKIF9+XaNs0Pqp5mZvOiUcDpz03yljem
2QpskOH9Xr2Y4Mgp5tgfx7/4ppm0/eewK66KALuBeZT0w76CcEkyOgXmxwr/T7uOoX7cxAtoXpSf
ungLtEZ9QZpwXlbyMa0MLVUDKu0ktGZlWG414v3KbppJW75WRvaUCpLKpoPASQMuk4x4vpCnJQwA
KLB0ucSNM4MbihW1nQXwl3+3QZHEn/SayLoD7OTRLba8UqFdeGWoTZ1oztm0d9SllPxmfxehw85A
PIhGoRjih7HKVScDITMJ7uBBHofIHoxV8pciZQ46ZXwoEaaCJYG7LVxbDKVgMsUVODrfhepmTsNB
Zbo7tClf58mBW5mCDS4pKg4/JsyZqa8ga1Q/6odJoiAlJ0Nhx0PuWb8qgVCVPhKBneQzxqtacudG
PBpIZZJ2WDxLV3jNmcXr+G4coKWDQTnrCsicFxWudE4kkZyhsdmZbVUn2Yor78lwR+3+9MtEPl6Z
FzFRVyzfnza02hTdEUZISajTHqmnVZe7e3mktd2/028sTYIXvevtXiIMNxIASyr7dhREIg69CpIi
FaCf/KNcPcDjPjQ/1relIJZAelinnoQL05N666sd48v5luI3aVkJnhvsj+VPJ2Mn/Vv1OI7Et29r
kyZBla4IiixHA49ZnAGN/9lYUNoqKfaeDNLUpSPvwgCE8EZz10vJPuM0c3fNFUoBzHONwKHQ2r0M
lHvalVYMMWzQBp+9GOXteu7KX94xrcuf/wZrP5zjBMiLCUpp65xm+GObWXqI0GqXOwm5d/2pBPPH
IPLv6NaGda4sC5HZrKx66wuDI0Yww1k3ET5Co3rubAXwQZlDiZhepunPV0ArU8apwXHdHgZh1uj5
DiTNkB4zeWj0HsscJQ57CXZKQc40/gT2NWziU4HQu1gvlt3hnlspwDrGsvVYgZ40GiTmRcDiahU0
mnMjtA5nOmDkcZ33Icq2OFgr80rydtfv7F49AsILnyQ5CW+YwLyCGt7SwnbSJqfnrb8limWFJdTk
ZZ7VKnpw+IvBdOD+IYWv7FWz46Br+1K0M3baTrXlO6dZa2D3qvgikoq+/43a3o2HzXA3Fl0u1dLu
Z+8ZxrcZHZxdpA0a0kvldOASneAH8gxUKOZFOb82vZ8fx5On1iXvutwot7CdKFBGhXVX83TtxbYJ
fiWANRxkIikVNiWlNW0NdDqwpr4AA+XZWaQZtGdhI1zJDbPRSfRUCy5tZV+aRQh3PhkFztkbSKV9
XqBqKs3GkaEuoVrBU6awTwoECSjc8lliIRMvvt6kdP/3DI/hoOvd37q5cDtDW0l9IuN+UViOZ8WN
fD29154sUM+ZmBV58lz3m3kc0m30V1BUCgNv5f7pgMNjKi2L9uQd2V7+WIRxQLQ5tji07qgbAJkj
irSyPXFEC0rNPmwQsDNdFHbiNcRKhP2rqftqH04MpMl7gsvQIr1QRCAgs5joCqkc075vAQkkb9mz
l+osdb4vSL96n9DziEWwVlDiQ3gB2yC7KlA8VLKfUCp3fhk9r7b8sah8+oI019HTMuqCH+ssMCVE
G8K231ugjJwiVXA1XbX2M2D2RM4UjtUeQm5Q3COscFfeQNzCwDvBsvJdnZThMXj+tLXAwlwoAk0L
vWRdG3Y0zuEgYB4Xat5khk/osUdguPUZ2kjsFd1ShxOiV4Ro51Z8t8b2WMvygD9oGHRMaj4gNApa
WAoGApc7ziQQgKp9jjhFoM22otyvfV1Y0ECnZM1OdvvBwJeFvR0Xg9PNUhjAiIsBRQpnxWcrXOCH
BOyCorZmmYwEo9tKtoazQxEB2I/MvqUbI2fF+YXOb18aAQb5mm38czo80LqwiHhfZiGSa24nkp8o
pFnwRCYpKoJVCbJRQtkwx9sJrD/9rhZvbW98XSPfwKDsfURFjvvoKqcPSxFP5CUC1gugCeHQwpZh
HxYodZPykKUQCqIx++mTk/OtYAKsQ3dJRG6MVBVE4jDLIZ6aZutcNgEqREoIz/y+WfH51Uak6TLN
DN10d49djS0LJhduyd06d/+Y8R52MdGmdB6hdVdH9X+PaFeELKc09r523tsCWJgo9/VtTUv0Fkwn
AP8XN42ma3jHE6/EuRd5gpYl1ImJfnmO+/Kb4YAnHww84kACJ5EcAM43Hd4tRtotkP5N+gvrSL0Q
POwuBxUcfRUjUdpgKucT8ooEMmkxd016OEILxbPzeZDxP/TsSCJ9fZi65laQS3K5dMPLL8wSsxFO
MC3EZQboy5izv/McTsjLcHhb1D4KHspdrpRXl5BdsdhUgHsbXpzd9rzttyk8qH7Q26K2np93XRv4
txdRZvHRuxaQ+5lwIQ+slZBuhSxqgbjZ0+HHVyBbueec2lCAq7Y3WJAkvp/pMLv5D5sjmE91Rgym
SoC11F8HA9155olHlPU0sIzM8mRRiTWfPEA1voT4sKQSHygyW3oxs65kyKlWxtYxbiAiLM5FP9tP
nzNKUhFwb9IlrTGSTuzkB3C3eipX9YHWi+inv00pEXkczLXQk/crmZ44VUBDGtG7RG4BaGCKetHX
Fklkc7WRid81zhSFbtVCXhmMopZXxtiumN661aMLOFDg6ZvWwFb3Y/2RNwIACWn3ZbWhLPVpQbCB
/7nfRcd1cls4N4R5YhkZEcyk9j9gEcbz2NW6YgHQxTwATMRrm8JDj3D1xNFMpszV8fovgcrAuauZ
RHP2Nu5OsyEj8VEnp/clpTXHKyBycIdCOj1WI4USYGBtYhoUcVSPIgYVdIO+/l+x/6gquoSoMibG
KufOfFMGB2nlX0nzVWPBZrxNqiGr8vupGHmsX7sLW5PYXV/7y5xVJ/Drs73Sg3pmR29+EZOikEnj
Hzr3Q5yNzWWQ/6/2+bNmHj6QZ2DF+4AKNmX5pEAWXrxjxBSrOjXqqShrsCBNilvvfj2QVYDG2sDa
iyiIbtXTX0Xj86Wl9a1EYbojZFzsQC8uCGUiVW3ofyv75ZRWXIO/s4gp8+LXTfuP1bNwPeRk7Yog
AZK64uQJRHE2f/8/JJPlVv33ikt00c4YmtFZs3D4MLWH/Xt2u36wCGZDmLrtpQbuqCBzLXodGMAo
jDGamrRPNa3o1EE8by6CChDOUeuu5fZBvzJ/vQ4bVdV8j4MkNBkgovdksBaLcXkkKSlF6RU2Wpde
lT1h25WK4qRdOs6ScFmTFQ+YT42jIE/2idriDMAVrt2UCxsAgXwxfOnbf3jV+MjIoeXKc5CqfMP2
us6JMcLsrctzRFWXSqNMPaobUJIwc61WYbuTR0ocYpARShbR0JRWk5TNNIxo8NYTQl4FNJQ4qG80
h9Js+SU4r4zf6mn0Ore6qz2HBI+aan5aEWZHwfhfVDtoBpEV1rAQhJKgD3VG8VFfF+mtnZsAVfLL
L76FeFtTW9HZb3dRqSnHmhQDb40e67l1yK595DSm7d7pvshkx8tCnN6F7dvZJ9PPG7QqmoQbqnZv
K7h1BisTce42fv/oeyCARQif4y920rquY9hieNMBbIPGM2C/Mbxp1Iks0BnQ99GITA5clrbUmwtL
SDa8eJVsSjOrZQ9KzovbxEruNCkKVu3wQf33a2k0cDInMmbeaq+FoJbpFQuuKp9cwe1ttjwmWp4/
PS4YcBB/r6HNsDlaG6zJMHE7Sodp04x8a5fFFMNw3BMpbb3b/k+2HIUPdnxmwaApnwx/ZUrQ4a/c
sryWo2n62RJxYNxlDnsOpNZQMefps2uwS2LzhO6JXhhxo0DE2DUe+5RUY8dKymzCuJbeIUAYDgng
BMLr/1Gesr0CAr76cNUEjbGayL95Ok8RL2leDrhU0NJeliHVGn6G9oY4d8TwwxLi8o/XhpDRB6yl
1lC3MB8SdpoK/dfBYJpRv93yDNwx9ypQMx1UTE3yqojS5Ao9Nv+h+2klMUQRjn8wWyM0NWPFTjI7
k6OowRpIdLEm7qja7k0xUyR9019xRdU/3KFv81Nol6iBVCkG21uibkVaWZZ0RIe1vbV//Y5YABfX
qibicX8Pd9SzSxnuZHoCJIqq4GHRby4e6bhfCXVg9N0UzVVvzLFGA4hev+86ZuaIDYL4nPNMQxDD
2wCxjVMCfYjNr18vFGFO0de0TekL8Q2bVi/rJtCOGnMxGweHQ/YWoI+ys6dX1BNUND1Zwshys5VD
ujqBdQWLlbVkLMtPs7vyS+982wow2CWkwBioZWU58/w/PKMxVZC7hsyBGOiY3T3/VqoIYLo4qVEs
4RUTAGLGA2qXO3XO0SMNCSaZJaMs7y7lIYVsZXLmfb5ki8BhXeO6fYITBNwH8Ys5jkTh7nRKShbK
LplMxey4IxuhroA5rre9/dDXpJgOK4txCTPFw2pqmAcIsLCP4A7fAn8MNliz73TjF3XwR48m1ZUX
V+v9YS8YTJiYCT4ySWWItPBVfFWjm+N+7EEi4o5HAt+1tlm4MZDQHVCk9q4D57+/St3y13lgCi2T
+BlXlpgaMPBs0+BDYn0rqOraZNf0tL2UG8RwHYwpNcNGfnnthZVyHu7N374QkLjkVe25YrbbUyhJ
Td4DGE7f32R4YN+cwZc4MJuntibl6+rzRWyp1xqQXfSWKj2/7r9V7d2TaFab0odj1thHzGqxJ5Yr
uRrQx6f+unas/AkGFJvafuomt4ElJ+mpkkI5kl0bayLa8UHXOi2dn8Ynj4WOpSv3/d7mDCXVPzdu
2E7UIrWnEweSkFq/Y+AOWX3Ogcz62bpKK/dIeB90rBO4Q5IIa9a50zCzYG25PM8DurvuEgsexIms
p7ch3MnX1rxfXzqPN27OgdFyHBteBCadxYUmEs3C/+PGRCgUvBTaUnbVFcxA249fxt/AKeDiaTJ+
KiRSXAl9EM13t0U/aeMNU/c5BK3WZGfh9uXpujcpzqglI9nzlVrvxLPhBw0VN5Zn2dx6EhXsAneT
ybuMeRVSq3qppFqjf2poUD/NEODMt6gY/ocBuRFL6w9qnTnrmkvxH2/Ak/wjbi+OF0/QFADolL3O
UbpVm2mxSIGiz+f9+5nGDVZ4f3jeYa47yWXeAMpEVDQFmcZLZYIj69EiT8Lr04mJQT9O8CNIkSBM
LYc+QZa4kLaQe3WdsuhNIG04oB/3sj0cYRM4EqnVOk5z0E+jmUFKJOI5fQ5tlBxDI1zC0x3rvVb+
D+jlZ2jnEBj+EwtEo1zjiZMwrI3v6/zI+fZxpWhAzSs01sJUBd6+P5qU8OPYq303IiZURuw2igGH
bqpk9XJpCQ8k58j9cl8qc0kuW/M4OriTrqQK9raoUK0SlVyPSCu/ZVciuVMDSoexxwN8hoFU/+iX
W+kmBXaGdROQNcJX9tLaiHT3TyFrxcWnq8+DdIhj4nz+3IEOqT40KoTV5NxuIok5He+2LZfKf0U/
Xlk/Hmb0hhUhG/4DVTsbfifxtxmuvoLq24/qdOyYQWAXPln9ym6wHfZrIM8AhwVVrkvuFv2BjAFp
tmsx0xiGFMN+IK2Zbqq3ErZ60Yd31fmAZjmdeVbgC+GYksSJ0rZH532OYlW8fE2mvdZuwvePV1wS
aEDlSbJLTR5rtr+opMrzEfUKzhx7uj4r002q7tui2EYT/1obn3Cz+qZyWRKgxF/ZPjrtZcfvuj3t
PKtV0qvCHZAbqyPCypGk09iQxC/IT8tpyy2GpbPO5T13MzlKI+9PqD/TI7w4DuDMaUXUKdqYvlup
YRr9hLz9joSghbKPvQ0r2tH0IvGelpmfeLW0SQH48aGqrns07D3EIN6N+plUmTpb8aYfMtYwK7md
rqwdM65+XP+iuU8a607wxrtcl8EQppJHjhsoydxXELarCVq9Es5oMx1FFC27VkVExbu7gjmuI08C
J2W31rSDdgPayTm3j0JUTd+VAmH7ctfJZsfV4TMJq54RYWDPm+xm7WoR+GiQfGFT0hous9WCeIO8
LxK0KiUxY0hvO1/Thzy7wn56ds3dYlCCt8tE0/68Q+uH22PFfmm6xkNl1vanU85IujKIGkhTcaup
f3lu02HtEnS3KV/1vH4D2K0phu2vuIn3HdaK8TWGRYM55vmtHxgAX1l01hVkE6lJoDfkacpY8eY8
iBUCnQnwI0ZmgKoxLt4KxVCpfLLjrg2KBjh3Tttd3rBsE2M+jCwKhdKXWU7lGizFZc2tw2jiJ2uI
5ysjOafrKp8Ux2exH65d9t1i45qxEF8MxwSvPW9H0roNj0PFh/s17hixHx7cEXeM0Cy7CTgSXy2p
Z554yKJThNyaagCGUVz3MSaDXXtdUFR4zIly1L+WQ6gJ+ok4tNg7YqXHxwSitFxCwmaeixvhH+Ek
GkBCJhcWMogMZtGl8WT9ZGY1yoDk8oIfNPGDsoTwJzMFFZykw4zSCa9OoBc0qZQp5nAMGokfwRBY
f5ASWw1XFWYvnbRsu8Do7gYKPhxKmHTWzank0zOYbaPVcgIGDQIjzy9ewCrVBoPkoFIeaicPQGC7
qUFrWaLKNv5H/pFzy87WyrGbdH6DZHTycrbyT4avxVgzAXgh9qd2rZK0rc6o/sl9Wvbzmk/j7z/9
cZLsaSH7ZPOcoaYMIN7F930EsFGoQHmJPq9sZxhkL3pQ82WQg9awUOQMkho7UpUhopYAgOM2mN2G
n3lQ9wJu2oBKvjzcQfgpuGkAXLSo0mYPGufzg/w2blZ/UtAI1Ue1pMRSPs+QSB//SWnGK1Ngwhdr
BmaWQUEfn+uaF0iYdgTQrarHt9zDrK81ldDL2+nFwHoXOwuEQGjS4+w+hyhYKhIoKPjDMQnzuwzZ
FdQTQyRnk+qomN+Z3fb4oeP4Vq7gwKsNQaQYvWYRRCZgBxddXl2hS19WbxNYUJP/5HwVAhaN7NVi
6ZmEdzy3Bi1+mb0kx7fVVsrFdN0bRlGX4Y8zT5tGxxZJevqnXFvC89mGfhu99Ybqee2HgQCaNVfu
eHK+bLa00yM+2AGqUJeullZjKSK19hIMw4WFimQbeBj4ggiU7xTp5XfcGtEIDlBm054CKQVZpCqV
hK9NYZDlFVtwQ63LHrvu8J1fSI7w768c13+88SJAQucekVAB3C/EugccgMYkOsuFotQVc/+iKT0a
JDyikOi4B4GLlfgzvEB0LggJEjMMCi4V/sHlWbRfFDsYKciKOM+DGHK8Dp5qTYL7OY3XWdfGB71r
aZllaFyNz4C8rUZJq34NISXzR7rcDqPusoJIlu2+Vl2+7H5NBFEFk0o4jPv6nphIAOav4+FYdcpz
5oD6zO+bBgKy2r9yxJ/IvcQ4sDYUENszmODu/cK1buiP26+YUx5VKvK+Mle7gVv/C2r1hlfJVfeH
dgc5p0DZgbDKuR7FG6ersRsS1eXI44EotDjw/FDJAX6fy9lU3Xs5Iewpr2Pi7uuoJIoc9EZtxj31
+1uKvk6UIbrEodCJcldjC+uQFq74K8Q43vJ/L1Y9lX+cjOKSCRBjJhi4dqSaQR3dnbqlwsXArqkI
UeDeNBwVnx8nzeZ/kKgAToAO3u3mwQow8PXEjLBGZUph7reSmgaCpuXXTWDFfy7XR6JauymPuyTr
URlBZbQUHq603o9IfJ5eQfrkT906WSiZD0DnNamUh8nCmoB4FpRHIm03cJbzs7u10wpGzb8vTw2u
N9AD4jE++IPgH00XgT3ZYSmEPBZzmDdsbqP/7YR36qZeT4TKKsclgeiXzl6aFPXzIOxwb/Br8FuF
gKylgCMVV65VPe2nkYGT5ZqRk851SSxVW6+DAqbOXf7wCcb7lbQ/bbEjlGrcRu5SrKTDaCHGhtmO
Elsv8ULnSZYBqn2tWPl4kzRaUE8TFTMc2NzDyxtgou5JOzoOlr7IpfBacG0NP57E9XwNaKkE/DdJ
z1f4NocXaUUL9e+Itjis659VF012Vm2GvP+HLjgQtnWqpCkB173T/KNWkI2ID/Bv9ovakkOOIztr
ov6LzzdBhvdQIqvGAKG8kzwb4MUGEmmeMjbPNYG1eVrKQRAfQmT258W2q5WuIhDCX7zABRFwQhDp
JCYlIMjRfVnlOdjN+RDlaG4DJMPP4M90xmZL7ocJHPV1zHvGBdDh05XF7B8eY+q+qeNpdrNEgXrs
vuaEMB6saqU5srIL16w8M7w/NsPPiwZ9QldLPIuJAD7E4OiVGgVNQKMRb+UkKSB6nhs1v7lzu6hV
r5o7D2FyH1/OJhVt8rCFoheXbUFBzX5ZUCUjZiLZ/8k66puve1TQgymhL/gRXMqkxgoWIufYVoK+
fSLqOEQ55wfT5f9HctTNK3IgWZA48bD4Ziw9yI+/ps7kmPm3vAP3IQCixpBAd1vfklKSmdo/nT9B
pRCfnyBwfOneVbuqRoyU1CaQ0Fi3GLdwvoPKXHx13kHccleSmkaTerGns5iysk2uhC4s+21ozbTT
9hsyZZ5+vFkub6FljPJLVxdxl+aMtNuRG8EOTkz044ZY3k86arFDZNhHJyRmf6b2gRcbG/VAr1/T
1WIKWDFbp7jh1t8M+nSapB3pa7sr0rd4FTmwO2mK6Y5qN6FqG6EmEpwZOSrLZtIqLdp/gGMbeUgX
UbgQp4Q+ag3aD/c6Xfh61hlRiQfaYwIGCDdnOgg19v0J9+i9Wnfhdx7qX0SjMyr328Jf3Rlls6Kw
TTabr8BP6Y5GB6QKk5OF3I3j0bRQYIXUq54ChKb30slVlpY8PstPGEWBXWVIn3k6Q6bjqNKZykA1
mM94w+648kDWed6ADl2NF/vz2yofpb72aDzutOdwFS/OvX70Q6qnIubTdZ+8KBghC0nK/+unBwfy
w6OUpB/D5zW3YyrIwnQbbdoQmHuPyDN+/o3v3P5XgzS3/yVd/xs18DR/tTFHmtEQXVlnnnw4D14A
iOKFI2cLwTbE8CohOrtn15L+xeupxZQ5T1ST1BBxIGGZMONf4Ue0aBPRNVTRYrrLSOwVL95ljrkF
Yl0/4aGeylyv2xlL9VJJu+rTs6kdL0ooUjcHyykTBulXw1ALRErY7PvEbLyRR2cQ0aHJsCsaaCjK
fL3Rf6sNVhFSAUvVRh0rznPavDjZFnYjYEpNtw5DS0qP0U4P9domhc38Ytimzzp9EsiKq8NnAaxR
Of7g1i2QAxwTCWYj+FDrtul0jUtC8o4VMK578TUtT0fHzfUkqF9pZq6n7tbqzlw/koXNufdfgJU5
3YxiegpNA1XK3eYfZWGWUGsETYErOlJf+l3lCllfO2zHvegw9eEC0L1sZ75COP70Owf2Ep9CRitp
BCCXpDt1uJe0hfMwWRgWb+7xCTRzbfchklXrRLYdxpz+zWgv6Xfq+CLBA9u3+AzleSdpRkN0yFgJ
4devflo/tLKIfrVn0c1c5hgIMGCBDRPwBMrGoJ/NLRGbfwIa8I3EJR5IOK5TGh6WcmKbUEcy5z9L
eUaNs+oPdzWMbJw/+sTuETqdzPV+qjcxsUlP/YSz4U/Sw1KyHetSzHujIeU/FPHS/IaRTWHT7toF
X+GwsJ/fs2KZ1b3b2s+jbH7XdDWQZDrTKJkzn8Nw0mmPdYnQMHyfm6YFFDfUI1mnaulhx/aD1taL
279Xy4Oh/SlqVOzNS/eAiT62NvXlhKFXKT/L4eHcr+joenzeXLxQsW9rKLhQ6skEp07nvvR1gNBq
GzvPN0eqJr2bYV+lfGtY/tTIbEmJQT5ZXi8XIiiH3bMJf6jhFRxIB8C29XeS4OsZlD7Uau8J9ZEx
NSBOdAI6Z7UmApSwJ6kSyHzJyxyGXtoZnyW+TWdVXl6jM7nf4la0GVBg/cQ/SEI+ldIBWikgGvo7
EtD4Kj5OtDXGemsyDfjkuyi9ARBi3pdMEBBZ1/KX9OJ2+Z2LbnDzhKzxbtfRBvxfJVErLZb0r6gT
OJRk5GyXaDHL6nPlblGwRpVu106dE18thmbV89AeFAQ1545Jnb9UAcI29a0NEuNjxvd9JByDfDPH
PnNJ1lqn2E64ulDwfWIaikEaPmSueBDrGppNw0c1LPkOiwgoOw6cF6iHbvkS5o/ne/rcEpBaix63
nnSJpos0RClysqCqVYujIc/wNAjqM7epQ0j51hHOmI3rWdtFO48eptEPYOtspUB4kPWkigPJqivL
7yx2aYNEOBD9ghAfCrMM6h4zy7HgSjHYKziqKYWLmKH4w+rrrYcBTswOt/SjFz264y82vRQofRw8
BRNfJICuPaCdj6efDj34gIFYgNIVlGXLK27vNvJMb8aOwispyLzD7rkLLdiqao3IJYktxUiU6BVV
UnMgYLzJcWCI2rPOQ/30lKKa7i/MqeIG9N2Mb3eyY0SvhqK15+lKZvBPoRjYOTKP3QOElq/TGdOh
2I5YNFpnYSN6FnpJDC6wCykD2uGoa2JKXZAgD6JA7VBZNcfkj13zNkg6WBMk2PSsVGlx6ay+L4Zb
mwbAvlySlVl6l2x9YVoGZK7Gh1Dh5kKzoi1H5l98tzh4chB/duPckuW/0hDg+O+J1g9OCWbQHYNc
fD5rJ5E5Ks3QeKf3tcDRg2o4hNIByfDDn4YDi6Q7HGkrRfcOp/HNzNoy6EFY3kootv3SLhx95HXN
IRz4Y+QOz/iff2wes9yfb1lcP6KfmTv27IEyV6F2MMl5iScqdU0m10ZxsGq+jVaOY9nokrhE9oCv
d09nryuVELUaY+xnC7R0JFtlMOcb5TbUzntUVxYojCgVylZJpqQPnqy67ugr98+W6G+DdAxc4PNi
B90QSkMFPTefV+myJ6VNcfGhHfeoN3f5C+kywteAq3S/GjNOicRaWcb3vpRNIv9wjlWrImk1CGFj
K6h2Co3nssif+TCZJdcKasHjIyxcJrETcecOsaltwcRiOBBNqMT1gxHkNXYFG60F2yr4t50DBJKd
Z/LiDFfkop1Zakv0ZRJEPMWHynyFpZieOyUu6AG/cXh1sO8F0jazhhoMhThb4WZ3G0YdtgBHvsd2
EgnroEpUj0IUpkk/FTnGYpimSa6OHIg56MrrVE6llZKphKdi5v7c6/gIPiynNtQXOkgswqkTJw+X
0zViTahh+CRkpeYEJGd750YjTbgQC6CecNkBEMiSwQPh2SasyxD8hVfFqc6E4k7dF5ZuhpWStUz5
GB+7HWoksXOWo8nLCkEQLp0Dx2fEVkjSnT8Zd8kTGurccENk65rhyjv3CR7e4RWpAnoN0T6RK8gU
sg8mL05JMU24jj1c+jdObZKZFuUBdLf4IKpKqzZCoFSXBGY/2Ihztl5hGEDtdIfJMATrTAHkik4D
bjMaYrSxzETHiFaOjUeyglWd4uFnoW94N2Gawfqo2e5RxJuMayqdhW7rAQ7eXgDoIGGJglO1lpeE
AvnTyfRI7LSoIhLbBtmuakJEfrNDE69yNK82nBMdSq6xefMUuOAExDMRnplLpcEG7Vmrx2fWjxXt
PgBrFWlSoCzhSdUj/ax/JkwA5KIgLra8TmGj/GnVzggWgHbXkeKG8Gas6j0i+3Eo9kZsLY9FoDgh
WUoJTBF+WXEFGQSAKpR+FAiFd+r3vvclxcnYepqOEAWuBcyDXuzF7tCtrezRQGkVShzrjIKePQ8f
QBvcz3Zpb1AuD7nqyk1pRAJXaBbHqLsA2TQAfd1M8OS5P9MS1i51a4Hftj/0cwNotYrfgxwDZKM1
7plaHroVaiWjR9iFrmHT1xqBBMurGPX0rALjSsJobVNpjiyC25lKpJW0CzJabPdfASLw80jXI6OB
O3rCdKoD+wg5Qh1JbrY/p8Ne8yVorReyGRyYZZJYz+TXQ5m8YzPYLMmU9Q3GOvrK6RNuGEFbXpek
s2+AnVXWj4cYuw8rEdQQxTd595BIoUv8JseOB6d/CSBoJ1IJSCjsKouG1H+1HXIqOqz1bjEldBUe
8Zt4QA3KHTmrhYiAqtbB7MNHKpHZPelSDqoSPHoPuOmf93Txb3XXAnDIdW3imSgGyfsKb1rUZNI8
5uVeADXEUDyAo56rDQdCBRrxkBvV4F/6sj1z8MkcE7zelILNgamDPe3FwJxruw10U5I/LpMqu3TD
HPjdT6pIA9+DrMC2Kq6kYSZfZtjoS3RjgrA+XXuuEFDqPIULkS1gTxTRxdQ1LB8QnM7pxZ6OYXV6
KODAcdmsK5tztljodE0g7pE05jgGKvarD2V/RbiD3M7O92n38j+na4kWNyhfhmd8zSGndCh2GIcl
2ihzNXWv/cepiWhFTGLJk0ZJNdY3Aa6FTyHAPEhj8G+YGjsQdkLosuIZ/unOGzUyPygHctlX3D60
Rm+ku+YINYOeDf9XSi+nUjqOIdI/K67JTPMIy5QRtqLXD5PQETYDxaFQc7I8kYaGHJDDdpDp2EWh
UGwZiasTtGI3Mubs3JKZ+l51JCar2K2Rus4oO2U6p3rEej1PJJurPUyJPa5qRNUC3JJQWwjf6r2r
gktWX6sMUB4j1HP+ugVco2Ht+WNI22ay5NmcJWkkIP6YCy9G9Qj1VO2z/liI4Xzpp6xj0IPCm6on
yUVMuG+HjBA9Wcpb18iIouYvs3Ks/zLp4dp5tIrNnJ1cloK75d4JygtfvfpPqisZwkv6wUQb+TbH
uyIPeYx70nZPvkcuhaVdpZd2zjyz3Z1SIfgV7GlVi/ZD1DQGbLmRA4htcxwgp/6qgW4gELHGUBLg
IFX8LWaDsZYuRAgYtE8/LQYvp2KUsMHcbEwp5eT0c69u8tghSwC+IlXxbPK4VNrnUZMEcrd2eQRP
wAAfr1lA8xlhRe24WPkXFRq5Msnv9FilVh1tUb5OHGobwhcZWuhh4MkyDr/6JfCZFX4HjNbm8/al
v/tW5ZkQrq3XtD7kG4bm5auO310P/cUz1eYvhJe8kuHf0ScZxKvQvcMKK0XspoQ8f22kcmnPhsjp
vpsIHrqWbKv/5Wrp6CX8GlcH9V9C+AEVi33cE9L+AUoT03ZrnnmTnPdT6waqOzlHZgQNI+Ke2NIb
yvZ73f2BBsVEwfXU3KmRsGXSnRcfy8drIgnMTbDZEIWrXR8lEIB7d1UvsKw6IcQKyMX48aVXmyjm
Ki+nTqvQ9MBrEUNOvoIshp9HictWVzxr7am0hBTzMp6BWZOqtTI/ZmeaqpNcsRqPXY6QRc81595n
ShsOKxaRCswA4rjhnaSiQtYlHDXaHA0Jseg0nAxNEiM+52D5sXYQ0nlVECWnIp6nrb05ez5NQojr
EQJjjjPEKlYiY23AaiY3b4jbYxLhQgj2Ly2FpfrmbXlK1E4eOoRHgj4QxT+6hLRiFCOPBEojwrg4
+r4u839+O86xB4trgjwtRSW1amyE2qIVY6IyKJcaBccveOVEPukqgA9KVK5n3jl0FUkXrsrMCYfi
MwhAIxBJI8Hnr4auPsJcCK+hV41ZZil/WvmPBrEK09ME/1X4VpjFck/PmPAb8JZ+iEdGqObgSRCV
fWfhoILeVw+SyjrahjQtzVXwJd5+75MPs/Nm/kEEAQ2mFATyKAQGNVuRUMV/aoRcTfcyIQe/YXR8
txg+J7A9Axp67lZfjgLoURgIDCcZWNCVmsBdo9AMmwRf+srnUnsdDhIPdoTKPZreeBfC9WYTV5ym
DKoz+beBXkBZQ++dYYtWCO72OiUxj0klKRSsUjxIsubPGwZWtgAnORKzJVmab9aHEfcSXtMSu2tj
T1JhPxFduxKhPajPjf6W/Oq1R6m5BCWsjfDjMBAvyN0MIZ8U6HRrsOIQEc49tHe8IMYAwmMhydoE
mmvoFDuYHXObhjRqm4jNLY1rkPjnB5skpiwWtA+d74VecqoNN2qpP6EX24ylkZ4Tkoiw1XVUZ3Dm
IqICqaDrlha8zRz4VuvkmxT37gqOmOI2o0QZfic78EdeNWiyyevn/xI40g9Nq06OGDawjX0sgF1y
9+axWRXoWZOjxXN/B1HY7gTPywVSc44yhru3yojLKlRgS14iyg+1x2BEs9rWo+28dJJ2Nyqn0u6v
c42kAoo+4wUDh5rzkzadYzydCZ0Kvjbhi+jScr5n+zanoa9P9hKxs02peywvMUx9sGDQvj3tHVFm
DuVBZTOa8Qiu3zs0v5gK3ULJVnA9401EwuMaCjQRz+Luhxbh1ShXeTmTT747Cnryvk+g38sWuVKL
nwcMHtr6KAGfRlvo7RpYH66N8jfW2m1YGicKcoFiFOP7ZBeH8xAvAG5KxWBqEt/zNBqX1ka2QW0W
BaTJc2/iTMKDW1daQwDJT5AYQBhrKfOdl/mUBGuXmw/WgltxUVq5/dRufNOqq/OM0uAMF+JlNLZE
iRmXIHr8IK4+BXQCq32GBDJwpbh/WKK8eDrb+UTqqmvzCfxgqkradjt4rQRsctArg9pY6cwuHw82
lfKtIffRiv4Kr1Ka71HinbcsHKYqTQ6iXKYIHZC5x9jbn9GGmOM8qt1nJGMtyXQZezKaAHv3ZI4O
ZSWZYkIULBJaL1CRhEf/5jXdLY9YL4b4wlIyoWqoMGSH962Ky0hN7jNdi1NNd48bqpSC+LYqVP/Q
EoETGjo7OR/FxizRim81wELiK3BeC0pwtgZc5Dq+yH61uv+DAvun20kkl3hrimhcKa+Yz/xqwEt9
HFtzMO8AkoAGUz84UHnEEtM5DuPKqyw9YTTimcXmgjFyBCqAgFLYRkaN8/v5YV6zOHEjfMKNRRKr
3fXJINxrZQA0DtQyI935FVeliv1hvu3N3MHjaicJ7ZU6eX3Sia9ZAkQhVetFtgClCEhOMOFVvtTN
wna2S3xRtj7kG/mVr27tFxXzFKG+qRrEFM6hy8pTXiUsbkmD9bNnP6fm3J/UyP/K4jh3a0WV1AjP
liCUey2pHH9/YLaduY+pv32TAc3Cd6HV+7FrfmsJIzLeo+VfAUowrRZhctOgsImZaLOeKvxQcnS9
UHm6xq0+t0NddIJKd9BO4Kh5KKMLcon15a6p7pKJrDWGhjyW37978aw8HXX64AOZhc2cZ4mLBQuf
xgPqy4zIxyfUe8hrIOLSDD8HzgEv1ssLGTkwgm9eCLFCXOvqqgPOluUIC7NQy2HdXgAuJ2jNZ+kw
wFfaJr504l/W583uncJoINuBZjlSBnfXrSg/fJeuUbu3LUVh2bUMJqkdjJ2O1gOpbbgAggZQTRFC
TBqSs2VaOD2g24Os9bLCnEUuyB+sh4h3MkvZxc2Czr/Ijh4RraufVBE13nQ2akfds3zwM7neS3Uq
6PF4fBx0ukAvACMNtBpQh3yWth2mCxlOkSt2/lFeDEYs0ubEnyQGIl4FEkyl2A0/l2ro5XFawJo9
NueP2IDjipWI+qfQ0hqFkbMxoT3qgBaL1v0NWXScHKoNjXUVvYpDpUgOeUd3m/3i9wfjVYOMgL63
c7nZw1a8UkVO6K3C036QT2C8v2sZslXi/TTs+/5nNNbMphYV2SwMekjonkVrxCPh7Pk5YGiRnJA+
jZZr1AsDcYrbAdqTHQm5zVYNRD+LLrggwvhABkMSm3xOWsm+OPTOSkzG1xandE/CdtJ3kQSPbS4N
5pwADGzsV/IRxClCdhfRPT5+uP+WK3Xuusr9M0Nn6l0fm3/h2g6BJlWrldC2CUKMMF4qJrsL+xtf
ltOms3YHD34ks1tYxvfP7D3Xyvn6lbHnZ3xP6Sr4AerYO4CvvJob6HAQ3Hh/mGCgFxK18PgikBNM
Y1TJ5oqBhyHfGrZbLuDHNKjnekYYqgtbiuyyMjyglK8DakM2drHrhWn94nyzD7EHpvI8hnDvs4+v
hvZEmE+NTghxPnHZfqNycS80aHnxhNJcqT1JMEzdPJfSlLVRsDVtqDOV7UJoUuw6agdhP6mOqqqK
Qo4MWZAjdxwL7Ic1w0mRqHADJSIjiavJWhWhYCYLDgNrYP8X/n5woWCVpOywpmRSQ5AUPu9VMGZW
5WXzb3A+zEQhhV2Y8Ckh+Vgfn3b3t1BE35lrbRqLWcT+JSlu9JSEreWOHpN5dLJAnPPyaAoGiYF/
kYW9vyKm5Sg/5zWgEld+nP4/OOhPZFc/Kl3yGA69yUVNSh1z4lgX96sEx8NVAYzHzUTK8r3lvI4i
+uG10hUp+r2ryTk1g9kidx99wqEbcWft9TWrClOz7lOis3+x9I6ZBRiw4fEnp3TMYK4Aj4kqycdz
TstLJeUSO9RHja9Ohti0T33Hmr+twqHRs4TiDOFYW09qTgzYJsNAKs/+BbJCWjqk6Ow+zgmeKFK4
1nJ9rrloJ98+jVtajnyEKYp+USZVHHk+x46HElUeYXg+zGKSKoRgb2w1FRhrWWlrxamQZNtJafOL
P4kHvPvTFogNY0lVf6DlHc+oAScXn0uwD52N2W5OeUTo4x2uptl/LucqudTeGxyXn+ZvVqDUPEMW
WyIa1zv84xGTarn41ct88CbIsWvfar3PfSV1EOIg5qCx+DhwSdsZVsKsEZJzJkXi3tmk1SmQiTpI
62sf09IoGXcY8gNm/DVKLwOP2TMK9rFkHij2PbG7wzPMs4s8zK+u3Z4lWTxqbNvMVgJ+XJb8GkLM
/Y/97cKtBfpIVvePqwzulVgPEAlE8xghtGz+4pqyg+uNdF1VFShey9EZ9exq/p0G2ysQpJfXqkAZ
vnPkSrVZIu+WfPEiYLdOg+G99p4WwNXeJ/4vOQD/Xyz+dT2q4HJGOu1yMS7YjOsI4Csz6n/ctJrY
pH6oMkjSMcri0WNrdr2E/PgYPffCHSjZ7DZWt5c4ZHC1pa90Lb3YMBYuuV2R7bEnuycHg/L3b442
3eGkKrkA5iqF5+bmVLQgEwHSEKVRyWsf4jZot3ypF/WKgTxBYH42sW4ZTbwS6Xq4dIgyfTOc0y6d
+5gWIyWua/JCqtq5aRaQMhqtV955luCj6vvBAvq6wEU8vGm+9q8xVdgHStppiRz2/elxlSyeZRUb
qTC7QwMr8MJppktBhfclv4d65875DGm15DBAX1t9GOoAIokiKaIOGEEXnqYufBzCfYqQz8ulAQ/w
s+tJ/QyFpwo++N0I31ePVRWTX1NB+rS5luqok469riu3s2f3ow0m3TuJNoqsoM/OgKAuWYN3IJ9C
tZ0IfocJX4xuQTp7KqW9cqQ3/PbuAyf9KzMA4Cpr8a3IVeDIgGPKz+AdNn0ljcNw7PY83PEevWcE
FGFxtVlP8RuckwFWBJcFSiGjlg27bLk9S6IBQVwYPjcH87t53Pj8Q+1O86DCENTUKlXbsr3uWRec
sTiaQ2Dw+9bGhjvANb7YnvHCWt88ziuzLcS/Icif6SHN6Hxo4vO5Y6N0GLmzJjnbJMZur8t4sa3s
KYhlqUFefxw5K4j66+/dVi/5PodQHxwfWbzDl6vDREagwFxToTXYkJ7cGdzunphbag3ge7eJ8KBC
sA3aD34qL/122PXZBaBwjGokSnoHfGSR1K9NtEBqdJY4fDdb6sswOMTfagxTU8LUpsKjFvbTCMnv
yv+f7inRwK9XzjW64E2tK3gD10gFad9Hux+zOQIPpa9JitfxcL4Y0q6eVcNtslP6QsZk4qxG+uBe
enZNdzmfYdu9OEkzltbpCks64N7YSILNjItB08yyPhRLTFKkJC0pcwVI3CsrUCt8RFl0ptq4vC+2
IIvEv63zGAqeUIWDL8t5XoN072Po3VGiwPVLbdkiUnP9WaD3q05/ui4WKZPfiDUZlWeaavOTwuux
Tzu8S9guBMP21atcIBOxMuiIwIbTYQ35aLBtwBUBTk5bIVkTWHkIxgEXpbrS75EZvmg/Sj2zxkPL
gbksqNZvW4NK7a/Q010Tx79QBR2G2mVF54O/sHHk1jFfzWWMw10P+pkX179djr0BgYGSlPMZIAI4
zh63pS8jQZOir1tQr4qSEef4+ldleMCmAmM/VV60Ah0dcEClLRJueEy/oklTFX8lRQtE2YQPONJ6
YReVkNbc7s/8I3mpi8EOso5Tq8gkmjC5y3kFtMnlytsVffzBN00a+AJyzwtaRiyJPfOQp4xGCa6T
eZO37NJrrRtV7H6sl64t/AZiNIxsubiSPILk8aEH2Ui+dY73zwt/qdDIk5ffZbVGf1yTmxNbewlT
k1gCrKVFqh0JQJrFSXfOnPnu75qFC3mADT8Q3CiNUlr0z3hHVzHHgC7r1ikW14/VZh+b3X9AaQ9K
G1MMby2l9mbV50okJ3TVVRKXdOEpo3BZ7ddkPK2LRYbMBbV8yO/OPhX0rzAOC/EVgHKBoy7nxKob
+MZ8JXVsdKZEVjKuEiwsfJKXtSwrMYra9zucjZEDvZlaA5z1LCempww/rigKgV3urnR/RA88WLoh
ELQPiVld1hZMwuzW8BHatbf5SLIK6lZOli+0NaWmwyNxU6jug5wlBIKyhlvkRdTxHK6qXSHXfNfT
Omg/9uoNiXJySxltPGdoH4iaRQ6Zk9tsUgYrk2Vu8CLE6L2kpprm3OgGxnBlG8k3xi+JL8FvFa12
/Rx/iPlwDCDv3XNoK1GlETnNjO3TngmVvT78cvWbkaJySs/t9BoAYFuO3kMTuYiiLCESIinTFLuK
P+gsu8WVHM1ey/x+/gN84mKH4AeIhtkvuFTfQFXR5HXpKB437BX9HrgyyaL7Zc24LZfmU/fXZAir
L6KdqsJrAMQepAvgIXE6aSok/lcCDmWZs3cQgLNyJAJK5LwRjzutWc54A3B6+RfZjxI87Kr1pCqN
O2TecCplIaoflGDnC729Z3Qn+8ak+X1OUHfhbJaEFwA0D1+b0LYAnUmuQgoSWz8pvnLLotQWgsqP
MI67XvWb9ljSSHguudNcYHl1dMkuwk5tWbTeNvaj3bQPREo/awd3l2+es2RUOvBXrraNfUb+6B5F
XfmJOkQ7lzWJwEJwyVhj59fkiRD/OGiEZBQcMsZ5yjGNXThNs72miUpJpCvyNWYG/HGyn23r9amn
SHasePlvRKnffBm8uRMB2FsMzHp652NXtgZeEv9n0JsAO40AlaeVb9ioEQ0mZPi8VQzkmutcGpx1
7aRrXrNsYBwpVgwJR8BdI3Fv7DiWBzNhLSVZ8pdLcRH9hGV0uolX8+3IA4VWVT69JjPEVFX1RkAF
Cee9VuXVAX533ck5V4qAQWcxR7jmQN/GAoQr2md87VGwTr5gK7LeIXFqyNk25uqYhOYJ5Z0YHwel
PADZWtiLbRXahgA7j29EyhnKmKxhHafsPO2eR0/0Lo9za2k2d5rLf51BGp0620Wg+20gRVg8eIuC
60g9w9wJuK5AoY9jp54OQl80EBTAjspYjeD0wXKcK2hg7UwH73lpWor4TSzd9Vycy6n34X6rltXW
C/EyTHWzvr9cSFDgNlrj4oGeVQQQIJbV2YV/slqhfdJBTNMJ8ceYA/aL1DpXo5D5bLoIfxFaIo5d
3TFIjDiI97sTZ/Q6CUmLtf0hAy4WlKYBeoV7tML4TlbSD1tFWONouTgqR3JIKvVtVu71aO6785bW
rWI0Y9/AL9acN8SwimtadFjo/7ogJvSdoc3wq5r2Z9JSWE3atoRb8DsV0ZnZnhVsEUZ90R+yXC4G
iiHOaTlQw/oyMXaqy1FgtVDfgmULep5p6iL7NBiYzFkM/anypTTTALNIcEnbbvQnOewc1X46htQx
p7S943mE+XRFrosYQu/+46KzOT7elvw8VxQmbHbNR5iVRIqDSk47glg236xXV0DCfuf1VGz7LsTr
i/me3lCH4yrSFpDm5T2R4cVW4lxsDZDUo3yPKJCesvKREAyrBQ0F3r74bK4U5sUc0F8iXClaLYWR
m7/uZT1IjfbjlZIQb3c3gLpwueLBywrzDP4irlWmQVYE4NahnGI4GnckaIv1riIKWeFe6d8vTMB+
CPqwi83wJdRy8D/urG0+xAdWamMXCd67FlH1B22Vx38vhaAjfQMWJ/GAeqJzviRjnxPgk0Ieto7T
f3fgDqJBqy78n/wSgMMyvxfkm0OipeuC1STfcCiFmisouIINNu7cmRPZYVjhCc4ritoRIFf6A/Q1
cAONc4fcB+sFwzZmekeyXTp+kCmwHboGUAqREbL1Dq7YE6q2TiF3kNBdVii7LvtccZnYrchoeMW0
qvc1a0oUPWwP025j0gRo+Uybx5IKUue9tCJsn7LArwASh24+qCXPbvh6/cGaKYPKZukmHFSR981B
MDVW+d5iUEXk5CH6vo207qhHwHrf41tp2BmZCm+znGsHH47mJ+qp45UNueP0cAV+bQJnUgIDk0z1
6u1FPNZa895m2jLU4Y8o5UN1dctgcZyXOfRJSBA8rFHWO99AsI2/fSVwt7YmYxoO4lDXtpt5muQz
LnASbYtYz5eKeGqwP7yOCJwT4pw+qIWYDTVrIzsGPt4QWqWpSO3IJaSIy/996vpthaQWJZ/IKJni
cY9OxxC/vnq9XBeGJSBzx8ePDu5w8jdEzygasLc9BKxH6XhunoeE3XjHVwzkFI6/e+vzsntaqTrJ
TCkCC1/iqQ0Vzq9KzQz71F1YoYVvYfrHlfWnEXecwoSJ90pSOIUhelIup8+XYOgr3Hy9DZITmoYq
2CASbdAxlA2oIUV0fKxqfNGJ3WaJQCMRQh/n905e9hiKHI/XwcT3xm36x0jBTTABxSsZ5TzgtOuL
AvoshMPRSYrwIeW8PcB9JF7EDJX4dotzSWEHETK+mDqP67HuejyJGmzl90D7vJmTJP/3S3Q8M7Wu
EF9yxBGf7pCh59WEvFLt3jedc5lphBGx3WKyJ9b8L9WxTPb8iwyPqRH/MDAmf0vL7hsIO60MUpmR
axXR/VYEEC5Q3qFXZWHzp0r/UyFcGwhge9J4G09HV0Clv4n2ZJwPx9XjrYK9KGEiJeiao4kilHvL
/Lp1ApGyZFryCWuuXL8ZSkJphrsJPhkZOSv+S1Io+w7HpzAUo05pX1gUKp9NEUMC3VdL13Ty0AZF
kt3h4pavFA6tPudZ8/i9GHuhIGOiICaZWWNR4Qm4EXsdae7kY2dhfv2+Gh3sYTT8I2v3su8b3raC
CdlExJqqNNGQaoBmLVlHPc7P14AxCJgj+9whpMjAde48D+HU3f155X3uC3sM7cnOuRpzIFk9SeL9
crmhH4J2IG5+SxWoa1nuJOpbKlpM2j2idnsDKQcOCuxnVnjD4QAWml0QwujbXs+bL06/0krFIMbL
kaZimh1JCnp2cz6bDo/OXSS9w3oBIEJwj2USNfBbSf0h9z4NrTJpAFIv+cdwctfj50VCBFfqOt/t
JagGjbkdJ9Nvs/lATS2upFQ2U8gWttMFc6JSh4RFSqwCcY/ZrJgQGAHLXsZqcEO+tyoO2fcrPFuL
aHrp5CXoPuqqCM6WHJDRhn4W2PKoiOc0X+AO674bXibPMheYzCOcElM9ejjcNFrw5ILYXn47qKGa
sLaUA76yhcgmt/B9HK0eT9y+5fSd1IXlHVy3sQMi+qpk6PUBsLbhwtB8KGWuvg3drGJImCnmISkS
vO84CSX5afTptNNIy6BearGGuy2Ew3dP9okKI06lGb+mHI4Wc205KPtpiWi9k8dUg2PzVdWBvXtG
eno0uwS3iSIto+wSlgfyCw9bGxIUvHu5ecbYOyapZqtqGBcrKtvTEniw2BeX34BEP+fttiSe95+v
H1/Uu2Uj+ptJKEaLeSMt66OuHdAOBjYIa0dpoxC4/NGWUC98ALXyIPqdIsm2KKAJBwjs3eM1vddh
fvtnsrpFJayoTC/Cc7NdRM9ctmjWOSrawONm60j+FiS7mwYycnqzO5X7LgtTYTwGrGR9KfHAU4aK
ORHqPQeAanCSm3H6y47oZYSLK1xSGlctgvzUXcV4y5LlgJGYQhivwJ+giLPfFiKRmZTUAVo+lx/V
zktw1L6MRjyy0s3Ry8/w0tZMbLgMrPDvawhdQSzDFeHa1YdNV99zEsc/S2ajN02Z1peK/8cYTTJF
Tv5KXK+a+ld+xulhQpnW2CwjVJxuasM0liKnsT/PNc1xE58XBPcRlNDouJRHfXedLup+zYec8S/F
NbRuH/LYSZryylxqzqAZapuQM5FvOJqeYYj52Ipbt8wOVlzCrQoPwelMpOq1ASE5tZnGtcTn59/x
S11vfjxWVLtySEdk/tBHoSra9VRTNyvFA/tXgCW+Y39Ytbh+DAmIEGWFWehxilLiVtWB+FXVN3AT
3HNkRo2+COHl0GVzpKkLyy6DXQmvljhpOWTt2d+LP4YnK85zLw5KdKvsFamYQSXbngRkxURNss5w
ermLre/UTg2WpOrHf+QcRmiGgcQlLJ1sc0C0CqQpKBXPInTFxoYx8wvc7TGLkew9B0I61u7K6WRW
5uh30PHZ37Wt8I86R6nAOqAXG0cMzLCnraGV5alK9Ce0xy1ldgreWpTMsMI2BJ37ATNQuy+3luOZ
WTZm3co+A4U0s99SZ60gxDVzasWL7fnExN0d47yrWItMBGJMcwNLOPSKcZ8RoOfFrZohWxB52KAg
ICVHcPuQ3I8FXNa4tATmcKRJ07GVOinidD3kvefpme1o4qNm/nhDmX0i/C8C06cpkuO0GAwCnkxQ
Bi6zKUbLOazyVD0kJ5/WSWWv4GJVLNkFksjWpBhIk11n01/hAx5/YtrmKgc+hTQsZNM2fueoxyiZ
cTelQ+qntwkjIY222Qp4fV5sn7Rh3+pBpT2Tenxmh3DAmcyQIUbZy82N2Joj7ZKlQ9QqE179N3HS
x8IA7yVDkrsonhsewbflTAdr1839OB4fZThWyc+WmOIa7UcOLgS13ESbj77Uo2kLEkSCiUdAX9Cx
cnrgbDwktlo2ag0EAdumoK5Szk3b1IpS9SIYodvySaApQYpaEZumv24XW1nBw/LCS4t664Hgov1a
a0OTn33r+XizCQ06yjQaTbFnLG00cMsnG1h+gb1fy4GXkmKjTRj5kE7vzhlHJunFp6lOCKmdDiP/
/8N7oHtS6ZUhJI092fu1lw6VG729OMUUNWpOoID2T17CPHRKnrhqepClB5AMsA2WZMDs+Y9Ca/Mg
k+Yk0p4TJ8N0V2Bb2MHrAzIkINUEDBXSCnCc6mECYzhFL/gjRaX8JXeW3u99EImlgzlLjZYvSu59
X7hSqPjRxE9sgee/QXmm1TEpsrAcHQFQcIwYTvO6s1bhDPaDLHgmA+8+YzeUDNEDRjTx71gbR4O/
zcHiiIJLeUxMeS1p0jgu/Y4iY2JqusvUxwS8ugWAE+HWVeXXBpS/JMN6WTc/kC6WiPnYeYg6i1YL
SBLQS0pjgBCNR1IFQkUdZCMRD1l9aD8iupwfny6P5IYCg6GBoGzVF3CvGKx3YHUEU9gQnrg7asCX
+UKrZR8oUq3XqLOgxG6HlblXcyUMDZ6mugaRt+fszTouxXsfE4w0cZe4nJTwVmSWjZWbhkPcaOel
4CdfUIDeUmNrnU90FMdvWmiTWJqKj0yFP5g6/dqBaLXcdQfC73qGsDdutSwwC8w0je6ko4i4CHtK
gUmgztOhk0goemhbmFSNwc1I3TAz52Z2ShS0+eQgmtgDMICpG8IT7Dr2ICOTgR7g3dfpRqWUfGzH
S8Shyk8r5tsCbA3bTj+G2HvR4JSW3aCmwEDzNxxY3qxGQ0zsWSa/J2Cf6p0a67LiqQYTYs41J2Tp
hNHGPaDi6y9OHid9hrk9NgZR81xOuSsoDZ0j/QNiana7D4GzJW6CHYEEpQwtJP2+j6HayysZlWdZ
6KulDcE9kiih8IhIVaUlyCIy6XjgErjnSXaNRACHCPDXI0mUChZYF4xH0YysNucYQQwBpSDp99UF
XyK8Srt3jQuBFHxZw8RK13Ry/9nxsI3NzUiwEa8tcccg3YOI9lTwyr3fBqFOFngOuk1pvxMgxPbU
CN0Co3h9wjG/2HTMldQAK5d0lcWCKaOhahG5WTl3W7EUu860rpGxtaZaEjq3PWKl4u45K5Jzhvfo
gPa+L/UUNF5uJwsXHIaLSnhgFEf8NV75wC63NtMMgrFmR4HBEdYXJgJed84PxySG2T/qWKJcirp3
/6fFv7jxEcaNtbvbs6rVoF3f68KeevdEEUN9rAy0X5HRM/c2Plkw88AbAT+rTLTNdmCT2yr0Vk74
Nf9RPJPom7J1RQCjN2T2tErMWMej5az42syNUbAV5VYrkyX10BCL1jzMj3aJNixMOg9bTglNBFw/
HHNdTSjsghYhBfbSuNfu6xH4kJO78oRrlRjKnROgGmxfYcb5aOnh9uI5Uf6hatwSGVStDa6LgOGe
bB/ILVBNPgtu7xbM/Ly3FIQEN+9GwQ9owAbdvor5m+X7K+Mzi46yeCRfYySziJPdNizh2tGSBtqO
QRPEGdxyPfdjM47xf/gKpdn75LAaaTPcVOBbuIh6S2creJ/geHHUSnmL9VXhKnkjXlIMOhGcKL9u
6N+wQ7CYBa/162OU5eUPDuYbzkrmUyidPIHBVDQ7RBoEpq1PBk0pYlkFBem6dOrvGocZkmxP93jI
GnphHAaoA3EwS+5uFEEGO/EInSRVjfAkSkvwGHh8DB2tpsUD0Kt8wsvLLFsofrO5xGDg//yUyR7G
6yFltcHOMR/SDB4VNok5nEnmnA2ZxdIdUiNt1j91Kc9VPTKk9OKRa9rj1kp5epKZwtmQt0jkukVM
KZyZieNSFFiK7Jup40LkZl04oPp31u5t/xfwd/JaOhTijyZbIoe7wWTWzPp+isyFszKLdjuaQfwp
SPN6Q/DMRnsAEoSF8r8ph8wi4aMf0vO9QVgDnI57zWxLCzuUkr6Y2MIerFobbPnGDYsrO/n37Ffv
vlpS4w4EXqKMLJLDK5BC6HrEA5VQSXyheu+hK1sZRl2zrwb6yPm1phhu3rpVt8fPMcPr5C74dp0w
3Gzn/90V67ue7AmojJXt8Cwz4W8M7U7A2Etc5ZV4AF23t3NPwf6qk7y1cak65XEjVXD30AV3kwzu
/oKlqwbsM9WKyn8cHU7ZxzbprBSxbvxrQi/AF0fRqbpsxMofRrWNhJMrqZTjp/YJ0U0WuoF6Xu1Y
B4LneYssBDfHNx74c1hKZxtF1k4I7q2QnouRk8hVqlj2B6l9TrrJcRFP+ZWIk4qi1UsynmBTFVSU
NM/Lu/K2RNlFRyKhw46Wi71R4ssNPYFQPhDaevP3RvzVlgTNo+YuuH/bgmEeJmtcQ9dfrp2+gXGO
mLDCMo3Gdo4RMLm524Ik693c0PbAaiw1bKhyUSaDetaGqzYhhZ1EOcGeoQiEhwmtpmnhFg+JbOtK
PUE52e8sQh+BvaPVuv26x6fgCGSn/agUu2RJdjKW/kMgqqm6jxVwHHTCFxL7B1m6UdLccJS8l0ng
UEbzY/wZfrZjWiKKp2uenHEsfHFp+t57YyV5tgxENZAlCumXCNePCU3bL+BaaIulWNA59HOENGXS
fHjM/8JwLkZcRcYlJeUF1to72Qb1HZ50XdcRJRNnJWfsnXF65g7S8z/8XKxVY9s1lJYu6clADyOL
Zp1uVzlItWnwbKsEDPO7w/FIGh1FtRtpUoOfwF9iXmnpdNjAhn5y8ccVyGFqf4CLe8+fQrJWraRk
IQFz9jPiH2r7AVhwXJ4xsmxm3wOadMPzVTDfT7QyJPZF5R/RNOoe0gTlpzRkFwlfmukKHAwH/wGr
iQo+1Xq9DPIcJws6XZ9KptBYgLohCyS9Bu1BiCq7pBcEGlY0SFzBrkzM+FrGZNlKOnCmh11DszOg
LeYDIPWC8AMdCj+jkLZHV0E5DdIpIBe0N306mw9Mpv5vg3RfiLetNKNLWKDWnzpCa/4+tvEtH3TK
5lB67MmfR9BGGFac2Nh2rLOwnUe+ae27nbboTFJj9NB4HPbbhDMXMswI4jQpE9Z5HL/owVFwniHP
drpcmdtp/iXXJ8op7D93J78M2Np3anzWVIe4863k2QqO3zR7jFb/9EGzSpWeV56zNmLj0IgnkTB0
7TIl4+0sOHd/467K80K7auq1DRfAKHzPuhACTOGOwVdGl2fW5Yx6m1qLgLb0V1R9fjbCac4eko5g
HT5GI8dipzEKtDOEPO3YDkuqAlqC/k7U4BUlY76fHMtjywDUQ5AkDxAH/YEYhZJD8tw5eGRlxr71
CBatQNCVulVfhBqY6aue7yZ16hjpFlKh8RGTZw/91PXIC3tn5G8NS1lEvlz+dZojhaigGtsj7NvM
MvknxwO/V8RwdhCwN2KG2eR0A/pvlKUL6v5LYKp/uZc7JK9M62DzRoMOYb2AcdIsmNXaN+o5NPX0
k8wtvdOU4lwn/roVVERR3rufTpK/cAEn0zialnYd828xiZtD1gsPwqA6mg2lEZcOYAxHIxTl3D8y
CXNZATEhKwoiQWs3+edctP+t06JY3d1ifQr83cr76QTEW0D/apRB6c/IpGIbjnaZAhFHqGD7naiD
mI2m3L6n/hjKHPOodk/l3Aghtnie9IiLWTtJJyqbCJPP9S9TVoy1T6RKeqlcSVWfVB4fQ6XJm5TJ
QjGTP0lwwY+woTE5yOlEV/rD+OjBrHpD1Km1GIvWd5MPLChYLpwRStS4LA7g/zIxRntYe7sMh+Mg
68Y9GO7D1Gcp8nglV1iCyUK0eDSsw2QX2qGq2Y3eAN6QwCiDXV6K5powMygXw4nyrdpVJZux5jfR
TSyVT1+0FtdL0iI265XlGOlLyWTiMgu44csk5KOYzP3MXTAjxDU0xPLscXc4X9QLK3TTNMWih8nM
AeXtPpApM54b/kEiI7f4D0gs7LxAfA3jm5rxKSf/kiHNS7QvYG5zyOSv874LeiMqgTFQs9iCO6Se
uuEzAGu94W5fnOQP1CrlYcmCi2nNwkfpJLJ0V9iziPuYZQziKfIXWtzzuZflJUvI1mFqS5JWz9GA
cE2sw8r6X1qcSkScf05t61TbSZ27snapafIDNEHCrDQp8Y0Re2xbjCqH1x9JAPpz0pFQ5UZPy9ED
WQq5yF0qB+uh2uvWYLxg6v/AB1QJTHu+yX7Jf/WPUBC/BEPoU8e5egO/2DmktikILb+MO3cNlDBE
5K79lgLDQyegSESKOZrSdqWVQc9bwemnsoOeC9QQfVzHtUp66/EFu5FR7iIF3eSFnPHCuHjX7Er0
DGDsSW3VO42g7EsFaPxtiFLu3lotWvCLSbC9eEJz+bRQCdYLgL40zYbIELpKlQMjwQXoWF1IOTyy
p0byaZiJii0jZ0zl3o17XftE7p+C5x2n3/ewwLY1HC4hrMDbUALxkY4DO8F0kTAyqadCrrZGDK8t
eqbrmJuxccovEF1sthK9bphoOz17GssUYVdEAn33cfEMMhsweM5coS6ypuz7pfLqLUpYltWagFod
nJv5lVVGxOLt72pIvneADVlGHwmJ/8JtfOXCPukEyb461Pzl7E498C+6KD8ndQ1jYYC9LFWCYVDV
GqPBEJOl33a9yOhIrDo1Z77Xomq4HUDyp2FmLJ1EllGYIg5AqRdfeAFwuvwzZ/AmQ24FDsminCdL
Wjav76h3BMp9VTB9luC/srj7H1gfWRxVyN/E586N925Gw4k93T4ikqsqanRtsKNJVS7XEPMUTgX3
nzrMiLz2TCD0RtVUipRkxMm7grctFAXZ2wsFdD3zG6o6F133H75SLfKjpJVjPImmUqMxFK/fV+6I
63lNoo1nx1L8zAazDaRapkMRvPfmQQf8z4oHF9XKb8RHjNqYDedouleinNehnYsJupoOeQh/MKbd
TwpQ7D1a+GpuIgXoPwFRcVnIfoJN5m13qIgqM87mgD+I5/Ny4sasORovdbjRMOTS3HvfIxGxKsHh
MM/ibxe/Nyuszw4bMKVaRfdgLnfnm475LDCrvaLHkWIo2SHbTCHSH5WWMheGCiQ8xDnqk6ayX706
KS3g4OrQ9AkLR4e1oxymMwYlinq7mx+h2yxSHqWOCQerkpPVQoVD0sKH9bbTuIh0R5I6IyyalcJu
saWnOzwjetyqV/jMqx46CC/MClg8lXOSv75Ue+RpX4egwIXLAxeSPVOpGEE9iWO8f8sJuiMLJsUP
oma6q6LFQx8INwsvol8At5tK3mugUwlYaLw1w+L0aG7IG01H2pD9VvbbKuwQNQhnqM03vUd2InvW
jaLgMBjmo7V3cY//K2ijC6SENp3NYquFDyukWacY9/mv8WZjgZv2ExMgN1a2vpd4ayRdZt1GFias
lp0WgurC8zjJ/sW6gUZflZ8W832wQ43BrRZjhUwqQKTCFMmnd9ZhI+HXJj/jn6gFrau/bTmuu7wZ
GN3D1T0JdSM5c+iZk+mQmp7rDW/51L+R5/g0LBlq+wwBP0GRrc3nw9yeBidPQoQQWJ0aJLsa6TuH
ZQyttZEAEBYTjmfp4yUlQGnihzI+lzwAevtt9rr/VPmu1Sfd6fZhlU1SMD+3F2UFL7vaHkpMq3vW
7FougoODsfqEWMiHAY7yvU3zLJZZCE/9pc5uwvQuClj6Un8B84ZoaLUfK8mIyIEecGjBMKSCPRdH
gI38KOpKVLJMuBW8Ej+gIEsxpw5WQeroalVnlgMIUKwet9lITHLzEatqhPPzcd7KwtaB/QdKGn8F
0g/0k0UJRyyEkYv+b/9u6ihbCXsHZMxUZkb0Y8qoz/XuLmbhl3+hnbC8ASGgA3eFyxdeYqgk18dh
oUy0YjeAYGXCB+YIHS4EGBq+rJAIR6cNM9v+wxKAgiNkqzuzrl58MPnQKQDZPWV28OQ9oaWF2S/Z
jD91fykBmj2zxokuCcpcKn1zzn1FPilxgGoxuAR8OYO9YGParkW1/bL4uaLUUuH8rF3CzcCfJ7th
lTdQQsCCJxs6Onplw3HEPqWPV1UvkbA9cbAFpzQ8ws/vgCkJTBLZFBpSpNzLx1NSsO7oasOPzRv8
80IWOHrfSAy7MEPlqMLHA2lqwAu5umwSnk83niEDJnRV0rloe1KpMIpuJZj0giM7g71SVGYwJdc6
Fk3OYXe6S+EXhyl9rpRb//mVEue/3SF9cDMFm1g2hPkE33s+6e3F/lOOS47IewsumDE6+i4KAdxZ
pm1aDeupyzC7xXuUCnCqhpRSsntDb9VSvCiaIJY1xXogw2FCE7atrJqoRfZORFMZOQDhLloiKDBk
OemUD5l3DuhNkTwnNA+j8dvkRlZDjc9a0dlYgCpRmpvD0thsXBZ4iZWnWGwlV/Xoy3i0Z/EEaza0
32oc2aBnd5cjUUGlMgUZcBux+RopMnaYXV51N66Gv5Z2fb7lT2YkfcP9vRz0fa1YHGoo0571Ia+L
tdfiK4t1jZHRkZO45AjJEpdATsEnsOwirMZ/PJ8KrX8DxTmIHlK7OLziRJR0pkBh8ss19r9bEJAb
j/VRDduY4t2TsT8nH2jYtLZWvmYby7STaAAidUdWNb3GRVNa5pax3n2Oc3NGttxn44EzlxKcJ1RO
5yVn1/sRiFTYeb4il/JHp+lygX9oOcQMp3534302z7uzAKbEdqqkjdQEf8YH8Z+2nDIwXQHUI87S
0hdEtX3jSL0Gn0mSjpDVxE9812bZoGNIKBYbknmq8Qv7RLYipfDTW3CZn1kqeFtlpahWSsYCwvla
nQS8IepUsriQZhu3zaeyK3D6qeSe8iBTExK874orvwhDNSZxPx80TqPwHYTEo86KhOHRAJrs3miy
nezJjnNyqqUSqESM1VttQiJorySi6peznJqb8xp0BC29zVrxo74Ot3l/768I/ronpR7/iMusxBbu
ql999m9wcxzWyjn007xLMe9RZnZzyIE3eYR18zB6QQ0SfSfjr3ZsEF/rT1MUL5d4KM+V+tFXgq2s
Fm+96mBrEn5hLVreEMtd60kzky3UTaA75+4COJYPphaGKELM1GxX+PyfYCth73efsc1sgjzUsWQV
fd+3OjDxq9W1WEMXjwcmoeRB6KaqL1zrLPtMy1Nc8rZ4KpmGMbbSIPpyN/I4HpWRjRfCfvLIiddA
GsDiP4bQXsP5G6YnP5QeBbnRbO2WxxBdL17u2szVr2cF9NFYgHnVmqG/xxno2HiYmQDUbe0ANai9
oS98sPqYNJisfQlV6qzhmwp4ewD6x4sWD+AWqWNlImokQ81ttTemuzvqmEFGerATh/+qzapiloI2
vS5iizzS6Rfwxq5azAAafMZhtDHSyVPrEyIlRXEM09/VVenzJwXsyZzizBwJSWfoqd25IVKmL+l0
FEUW7ieqqLiyHenOhQ5elsco9L4AhYlnBLJVaTddyzyODbdDPEiRJrz12YLcvtU7Jax6GUZl038z
eKKYUp0GiZ8PfX9SSol68IMJ879BLu4fDxymP+P5G77tQQZZFNOyqRIauuYPSKdf8VdkIREVCFE7
VpT4Z7tGfaDXqibgMAUrnaTq7/B3Y1KVTR333Fp1+c0jxkiyt6er96Q7A8jGLBxEsEYzUPq7dEQI
aAadAS/8epbto0UP2GT00yqqvIu8MIUqTX+P2OMdKr/lL9DO5P+OkSwzbRhklCT9pAiMAILtiG5l
orS/WtvBYzA+EOlHiJNBAK/dPjLpRaEUwxj8HHhWejjeZPVmbFyxffesC5ekrCqBYs5659rrNjGU
e6QeZCElVu6Pi/RaVIf+hnpXhl1KZ4AwYrVBf/opJXacBZ6REEbCIB02/Qk22ShBRPQZVwCs9X5a
AkbmiCFFbyn8XZt/5Wo6+pJhChT+oLXAE+x34uOhhWcdrX/Di1Iz3jV8y3iBGbqKxCJChhYfXWkg
u8KvJDJedaJ8QOQ6QBSuXIMF+tCzgqzvaWfGROfMk4uYV70hLJOGMM+Y6x1WRi84qZF2YNaxTtKq
+dJqQQhOUR1Ld4NQZJ7z3vVkNIepmRtoR6K2ytu0n/pUyALMmhHf1Orpt3sDyCHgctm/r7Z0QrlA
UHk3CKuzOcJf976O3C0IS6RFQngNfcXrKaObbQXjOpEdLjkKEwUDzulbc+D6MrA35gOSMIizlAZt
fmjb8ajLh1KloZHQ/HE4+X1DtVbwp19QRGCFZblaOb9tP3lmbKjY4UbbMdvkVycdqhq3VbWRUEK4
domUs356dPMQwHbJp8UImu2VUkuPmqc7YEDyCJA9wpYQsJ9F7yoIyZNd47ICc7ukG3bGqWh8y/fU
m6M3vXgoZS1qCDGWmUAazwayh4oWQrsjuP/Md4FVXgrsiTuz1P6ipm5M/4wWySKRF8JocuFJykJy
wv76X+tGK1dmFXnky5h3Qt9aWIWcRgvdxzc3vMKxP7AGT/mZVhsUNa0Z6YVlqu3s5tf5Ag1s5Lq2
BWk2xskL0hu3pTwey+A+KNmQy293k/sb9Vug9hZZLXPApTuLFPzrSP42tk5IzKsoC5l+ux9nKiu7
CWT0VfAGJUW1BgbCYAoj/AR1PaPJh8oZzSII7yz9xVX54cDzjnINsWc84b1DmXwwcTh3f+6ZDoEa
OsRNCvttTbjD1GEQNMcqVafdq24pTX1a7ViZUWauLFe7WG7Mx01RGgsdCJhD6zhEIRmumaAcKuM2
x4jzef7fYtrDfnGcfP5iwkRb2twcTLx8hUICJfSd1leI+io1KRqcIT6cUmgvpDHVDHsB+nfjtkTO
bWlV+zfgphX/VeoZjVwRESMRKMlYjmMrAiydGdtyFYaeELrSiU1GlJ1GKVPShqaIVLoMV+eTnIoQ
lc3rLNs8cPyw2zjtgjA+LUH8z8JNnexRwP3CvoyG9wCgJY2DHo/R74PjwfJSFf1a2N/kzHQ1NaFX
n4OcpN3hmALIHPZttfXt5oA3ptPy4Xux62ldGUL9tYdL76QNFct1Q6ZD/EkmLjBW8aiI9e3Mz7YP
1+yWmUlxSIEYzmZhIMxxXTxFkm+IizZMR4k5goop3g9vw+e+vZBOd+yXUWlCWvOD2gnAhOD3+Vlj
Iz1W2lSZwIJuNvlVqsqJaviPY6K1KQHUuxf7NawhD8b9Vg4rNdsHeWV0o2mMkvaz2kGQ4rxFwUjO
7vZgBw8CeaXEsE1Kuzvyq6acKI2U92jpt6IjrLaJ0W2kFZrdmfeNcrnSRrEAlbiLYlKBKFmflRm0
bUlNmy7F58jy8CnGUF/Pl+WGOL6PAelv+RLHhIQ032XrIh5F8EEKIpqmYgkMCSbmRqsSZHaRO5mV
I4uJllHSxk2+wXXCehK3iVaaaad83MvaprI24sJDWWAuF21lgcce1J3WFJT142VxO341nvNKWxF9
pQPlWcqoq/WeQeVBSw+2XIBhi/y+w5sgpMk4m6Qk3cxgH06b7EP3ipMxPwxOBfLozRVJvUyFsQVa
2CX3v0QZUtws9xDtItlqG26Y4gxOR/xbxmBS9gfAf7cIqwSIsxPLyQBWWiHza6C7K2RZxCSvLCS7
HjusTio1uGUy6cDT6hIPYCRvdLruLXZXVTeLMIrI+GuYZTezM0IhZcA/KXhAymNfpGJeDe5Gs3ob
NkA7zUrSJkf4/NMf4LcEfi7AeIPx6jZ+KfKoyfnsls8XJABYx1niNBSePYVHStzoiE5yvrllRV3i
6rmhLHjnGMMm3hPCo8yP0Sa0oHRQW4Vhyowbdx/dI+lqitI9TIhFblBc1chWAH+hbJsldn1MwREN
tfl5CxnrW9cF3AXL0UQottaflsdBKhoFUveB1fi+GD+5qorulawHui0JtCs9j8MqnPpgIIyaXRaz
TZooZoki058unVGwNTgjlzzo4kwZ5h4L7lvWTg/lwBX6fCBYN8oBl16/V7zRF2/vJryOhzCyEZMc
jqtX0WEvhhMB1WR8B1gUJbCKCBJyKaBHxWc/y6vb5MAu5y6Sdxk6cn5svXeKIDMqnlnq/dR+25dM
S2W+2tZcT9pn8TVLw0QimaGbbq2wspeM7HONcg8c1CO5GkmF/KFZFgOq53fdThVd6PkXbheLKZqD
DJ62GjVfvlOIcZEcFjD0Lkh7htPhAAqtOpwWGe+mDoxiQYf2Z9Wyy+8MPBbh/FTnp5dLOOXPLNvo
YDasCW434dJnA+GcBUn4G+E+3zgLVSljCqmrDyjxMjBduw60i1Gd5mYHyYGP444STD6AC3J64rIS
oFyXn9/EAUMBfEnQko2TOPcvrMjWLA0PoyARoWi+AI8WhnsU/fq1E5vSB10cuc9FPsU6IzoV5P2s
2CVfMkn23BCyTrwjfsU1PDIfggvbMO++55dhOlbux7t4b15uP9qujESSwbhxuOPVwltvb+6VycjL
XuwPjsDbPKCy/BerNJ8AhIODLZ4N8a+AI+0uOGJITQ1w4o5cDpMJFS3gkH8US8vpRPsYpiTyaSea
ZSzb54/z47xKs7e9yKBc385WNQsXIfhSoZTjdGcRsOfLabszCGoIUaRhl7A7TwRO4WQQT8WcVNVL
uFWHvAtG3w7nyS685BLRT8Am1Jw7ICRn0dyhQSuG3dua4AAuCt6PH7Bwr0HZdNIoYgBhl13zDhGe
wL5pXVRN5ka7qAy9izr+AaY15NWzB2hFAFrFshnpBSRLOJHtmlY375/pVFI+NxYIOh9/fBCEuSyS
EuaenunnDPb35RD/jr86H58UmwQBJFWcKGbQ6OozYfj3RmtEIg2Tq2s1aYBlvQ9bkUvhqWQ0JFMD
8xrl3HI8YVYdf6vvVATYnix4aK1tfiNll5C32FZ1U7AnhqKqeB5YpHRt1DNGpOBlXmZmlvJHh0xN
jAxAcjE9oQri/waoY1oXg+qNCOM/ZzRwtliVpspYWr7y1RuEBMDCZJAkUJeQwsg+zF/kkLJeiMHQ
R4wlWvgic71icJj/P0mrEYThsHSD0ZT40Ue0otuwRK3NK7dxEjMXvVEerq0szoEpUl46+K2dq4x1
tKvxNTytpFzijtim2oIH0gP5UdgrS3PI4v0qqjAyBROOIaLOLYEOTdMu6nS8nR0yMFQRkHSgMsMV
waHUMCm+NkjfNFBMfb32Cni8QE2Vwx/NBrmUsINOktQyKRrRlOnR8zzEjzxbwe2iIAygbZ6GE4Gp
d/g+hqiKdkYGKF02ZgaJIOLynPURTGETMPdHZJSCabc+UXtATfPVb46vnvBmSgp3cBaXrPe9xGrt
BTsKJhYieXz5fGx5VeUpfanBOUOxeNr1Id9mEsoY0uy3C5p1dj2FSG+yU/5f9EgceXef3xhSOI2W
NR3PQJKWknpQZ+gJFdA7qhYqJAjlN1yJnudHYSQE7SMHLnEiAyaeqQiXD1EwhRpTdD6JZ/0h1b3I
tR431aCPFor+Hl+Gq1w8kym3aQNFnwA25tF/9kUe52aYUGxleCv/w6j0FAgo/nNUOYozFVx0hHjZ
EFMEboEKa4IAURX7FEPpr3A77U65rDgAShdi2gxqfCB4CKINBVZi7uPyG+hXXsbM3V+wrokNciVg
bOT/IFh/Pj/u+3zY4AE+jDjjYdEZaDuVn2nqPFPdufphM/9HKu/0icxZUxiRUPObGa9VRGVBTvsU
4tdSct7YLeZ+pTgYzPcZ+WAXqjzHYpRnFbi7KK1G9qma5I1hFtFSTEQOrio+lnb+k8LpBsiR0dwc
miiSIC4m3h1K2OuBLcJyFGbaF2WCzNFQ0mtMwpFUr7dhS69Ywo+Qkw6sZRFl++2S1ijkzKgmqkcO
WemoJDLSFk1dlctDLY0y/IDVvk8ppQCLSYzJcHSfmMkFb6HVVaJqmFH09NLA41vgEVYDJouvmtmt
ooJMQ7GWxdw9/qbDazeaGneKIvxSX3IviN+oRXrNrYIRVhq06rhXKTG8Nc5NUDqmuKvXJIcQoi8h
MxUKCSIymNEuvTie0vR0AF263wOI+gqmctfL12FfnYrWJHGGHsm/yaxjIChgS0j5ZyIcXURe2yIq
+I/rEKVvBT4glG41JPZuetyPC2leHh+xQ4+iIP5ySxFGwjtgCpdS3jrlfdgesoDuHiROUyj76g9o
zf3cKiVx2eBwi2h0Jy6RX3Vu9wdcoR4gD1ajGsVeYECDYkEaZjWkN51HfFTZA/s9j7xnwJ0ttgx3
FX7tq0ZOyBLJUQFLT1W8Ig/7KNRj/TXqrerGV6BLeZ8mURC3WUeg8Zr45rhrgirNFBf7l9pFnEQF
3Q5bAE/148z0RybqeO/z2T/+YtAml/tnRMLq2YTVtnOXgfqFcJt4ArNBw8NVZBH+sLeTRZL958So
ygAjBsOQp2M/0JxlINq7l1EHIA1o6arpLxa1jZPtGIhWewvBeUS3pw5VFshkWxFYX7EgWuZplqWo
WU3yqw1aHdbbEBi0fWvOndErRsCIYmt13R6CQ9NFqhpG+1itn4Osls3kzlN5W6hkuWrsEDYbrPfZ
I3w0p/EoQPCNeD4OXtdS/uyWlOY9DImiymHSEhM11sz9+G1KF32NkFrKn2WzKxuPBW1Ugyx3ty4Y
tNEP7ome1T767zHkcACeEgYeUSHyzL4qjUjECpqOvMCDLmEScGloCITJ3FXAwiWBDSfcWKEUwQzJ
5WRVSlmZgAtcV5UO4OW//Qb3B9nVfXIyzj9Gf1anbU/Y4iF7cU/p84i+ZoVwR3alWu5XlqyV96JP
9RsuKBQ5UVJ8bZEcfyxPTY2VxcJBvw5CPc/K1Acd7lcNY21+3zo5Po4NTMcO6zRFe1y/Uu2anC87
fRUnXfkUB+5R0w+8uJhKZvV8amGCrqc89AMMsL25OUT4MEhNMB/z14zYfUTNXFqmKRfAhMJ4PNG/
81saigHajPsIK5oQhOHC6KMKtnPti0h8JB5JRXpI6YRVJNGcBOg278/YGDQ0YfchJ46U8+LDu41h
tMtn+CX56tmBMQ07c4eUCl5cO1znTSGLTaLlM/jp+VnhVdGC2O7/h5TaqMDMsqpTcblbNEsBpemw
QSGr29g7ofGFpN2lF5NklSo6G3UO7pBfttY8hatWBZjiIE4s+Fu9/FATGRIYRrxtqXcj5YLkZVeD
tvatIMV222m3jx1eM7uQsgkWjAWxNQnW7JvOi5p4fbH2BfVb4fZpsOlzW+HzsARlF5HfchPbU4aw
/GPsicjHvS3itvy64+txPDBvPKNHoDVQvkrjX84J8NwAxkLvjBpLq5uBg8AttssXSzGjlTqH4UvS
/eSqpE6DLCxkS3kQF3SoagUdt1RS2dmD1vLhHvyW8Wn8vgVtAYj0/U2R52XCvOmQMvGx7W1Fbjdg
8Te5rj4nYZjR52ERp/nDV9cAExfr/LO9Nn3quP72vyarsSu2O/UMDwWYEXxka6jlYEYaukwlTKCw
bQEs4HZmiPYoobfTVNtsbsaPQRfPvW7HfT+Bk2Q1C9kkCxlEw7W+61OUQR7gV/ZT/VyBZ9C+Qpjb
PmZco8hu2jrJDjf3FU9Ygo0t92DOx72Lx2fsqKtrD0Qdh1RRNUPJeMZ+Fpb8TmZEaTac6oWLUxip
mPeRiwuFKsglXsxzEvBdPchlFrAQxNRsgHWC9NIhBIMaJ6shko7CLswc0IHJUkCGWSGIgT60jxYm
TEFaFz4gsOeNGiKK+xFFRhyadyG9P6GrxMh3IUOr1TeGZy9NAxFPNEoeOsSrd2OTS/xnfXPtFLbQ
t5lvgbb38chE9mQrQArLdEtQvfDBTZgLEqb4PqBYo9VQwJoz1gvQU9mPNV2gv6bH8soLjtEz4gik
B72xjaxXVd6oiwjZyo802vMgk8lr4oBIBRzuMylzsv6fstmSNzrYyRMdmianyV79DFZuqS9oUE8D
ihf0T7KEfZgDQvzuSxVAMJu0QYD1/2nF6hcX8AkgpJPd4tasPyMHxoSIMzvGotYEHt2XFB87RBjj
0AUCCm06PeMr+dT9K39UXjxURkyVpBfzZGduKLrqBc6cexkJUmzZsznakbUQ5JlkyZJIndZFEBOp
wcJm1Akvvmf9xQpvlkKeJFFATJXHSLtFd4jxdFd+RXXh7FTCsYs7JOPZKFDe/pZwbQP2sqx2Gk9t
VQJhiQBH1w1CXljG3x4GaW3oaYU7lR32hhDCFIxD1GQcM5NZQWRTq94mkbr69Im+LISWAvU7Ujkc
U8p6LlgufleIJT4B5VYQzux5bQRq6GPotNINY8QaQtBJfED/fg7xp8Pls5VXCGVxk+FQ4ql4k1yL
votTw5oIoikf3LfOerhEqwv7vLlxW0ZMx5y+zYONAUTtNYCwUFdVUihiNaWMMP5YCmUxQafMoBgi
pwRz0LEtLgdmW+Tv8fvnP19XXtmGtK6QTd4u7HxhDm35L76lsQ6J75ZtnQN0sCp4hrh8vO6bRvHE
Fw3+hJJq1RdQwOpcuw08eioeGCkObR2NuSvNBpVHRL7VIxjKFEl3xN6kdJm1ampEIJcxta3MlbRJ
r4BqtxFpXAtH/OaGDfwgfBROKzAePan0ysdJmmCaTsBq9NpThQNieBLW0sW5CDd1i0Q0DNgecn0x
mLKx4UA0xwjuWVI8Xn7+hiIgy3E5F6wCEyK4D0XP7QRq1KwzJ5sHsffKAzxriiuFTpFxIFUNdeIP
jqeTUWHqCmlHXjbb4Z+oItUM+nIqOedjWsfZeRPRdgpFZyg7U0/VERPWTdYwSVuuvhQPs8uTydkt
ctHF5XbuXlViLJGk53CZTrY3SxYFAJ5oYbKLkihIXFxwpcfKvc0RdrfOzRmhatZE75WC+KErfJOs
II4MjnA82pZ/HtF9FCimGrN3FVK7K7xbnYw6pBxGdf7+615dGQn/EAtZx9H0uE5fB+8EvuJN/QzW
xXZMWZ6ZMmQITZM6k9JB5j6Kp1VX5kKQnrXZ/cwoLlnMzoifsLNoZaas7KuF1nBGyCxZN4kGbqbR
1QH1ouq2bHTsTuVHiTggYFelsRZutYbWiKXR42HwMhAb087CcLPhkMzBCKZRZU2DAFNQlbO5TKaQ
sGQYiYmi3zML63ufSMD4umHjBGTpwqA8fbGpnzlRR4twhfVm6b/+rDvvla8J1SJE3lACq7c0JxMS
DTvR8+mcuxSJWtBFsEf7yzlTHr+wKC0w+HnrGrcALmnpB7yfrvA8685g0kBzItEUG36YnYmHq5H7
QxVoHZCC6wDp+TTd4lB337PJ49Z43ks37yVquBpjlX6kIytF60xLpEFBIhHqAa3cI9WzRb9+qxJu
EOUBYNaU44K1OfpecVF0BIQzj1M37Mdm3Sv6LKQ5xQkDzJptE6+wxz3r/Hcp5Gk07plHLkyk8QI1
z+8mh+G4qkhdmO8W9HdDchu1H3E7/77teeRKlw89Bf+hQ4TZgYHsETpp2eIh//9Dugp7DzV1KHhH
JunIuoHZBqlGJVcUFlys4DXQhy38Q6cw+nfxafLM8L4geS+86vbNRO4guaW9en9UHOgkMzkb3bYQ
g67wIszsCbeIstgyjSz+zMlCIbGYUJxOSsDkL6S/xpKTVdk+SPaA7QgGdj+KAJZ2ojE/MvMZ2S6l
2YSfbQflCQrrL03YqWu0q6olZJ9/JUrG7MAutC3JEo4RMajScKvsW1L/BHmQYBPvtOqHbemk3e1m
SFOpzrBsXyuSeLUY2IQsNhj4NyyL7I5TRkX6s/erPxlTyiurDZ6blSjOhSTGqpQVvxhIte0sHWnb
26QE1OmVMpZmzuAGnlxSUZLHOCiddZKz7MQ7UEXg3bdwNbsJcTUbkaOyRvidWd33H+nboWKLQzXN
WZsxbnkyGi/a3w5TBnBrDu7F3vsnvzvZie2qgOu9FUumLpjkWSnLCCIFa8AfxvChOgN20MzrNQTM
x5e8qO331xrbCMJQuK/1UD8jklgn2mViZ4H2yrFT/I7er/iftRYzqmcKm1SL/9r/8sJmIdOIIe0m
2YF4XdPU2GVx398FlQerKJPmnIlV4+HPmepw93hmeFR9Ma8WrDVw4ojRp8+xRVFHZGWQi+VWi1HE
BwKEBJNFgN7Q+vqq+wsZHxmMZJkfPUQQTTqczB0Af+jVuAY7MwhApPKs8Yr/pLZKxfZIZSgTG4Qp
w2x7x3ahm7G4aWyUhjAJ+RAUvi2Z65cmIHJ2VhrGM3gl9B9KEjacbSoYTmtezSJYN2k3XMH2gv2x
ldS/WGc08yLfyW2OK+IC4j50YfReYeq3hUY2BGU1JyAq8Sz3CF713ydM+p5bB0m2V0mAd6uqEd73
rapuNBKWofpdtunG3m/dUf4mPHo881HVm2ddThvVcPFZ2MLsVR2fQk3FHhtVcpFEPOLf/NgNI5xS
AfTkZ7uYCSmB/qcdrV6/OXwDTJandTY2pf+kFnIIS0gKdo8hFO3e/m1psogqBfJln9z+hcSNPEt/
fhWLhHMPAqCfnDDJRS0LCTHFie+cXimdbhlzKMoCblZPAbaYdtohXQq0oGvxjTU7+dASWBHeyr+l
1TylVYWuwReSMNaMuwRVQWUk1iMBcmKrezJWhgZj1ABN3DT6YJ2xNOIfbOMymMa5greOMOEbnqsJ
A9FPZWTzXC4x+QLVd80jFK5AdD8F/paox2ni9dwCzYOfhKAtLl60b4PilJtxjGVp4E78vKJmw7/I
rqpO1jzIa3yD9qxnoVEliXMe+MqwrTyEE7N53URy+5e9M1rpue6R0DCFuwsN2IXWVlWvlMISx6fe
I+rZYeNJuw7PhPIDVJZvstERqMlIlQf1c2uRE+dlYOcLmUwMZ9U1dHUyc8bHLJmwWnljFnskOT+P
G545841XFLzCmR2ESnlSaBVziy3YNjvBsLwNMFWBTJN15qTFz0xiPZzucQN3AsDiPjAmKLNCMXMH
YWZVptpp31dmnQjIPIjUNfXS+rD7FPV7Oq/pZ0DQo40oZv9F9J5OYup9kbbnUwpD1boOji7/eVu4
rFgd2v9aaYTgpNiZk7BIN2g505KnVmpfG54wY7dy8CK5+J8wGNNTxhEnF3uYD+eJ8kE2IOLxmuZm
0wrrGHkBTBBIAVWGljOZ67c3FrBDYUCyY+8sNrSNwGamd0+W71JflXUE2Mbfjuzqy6YlYvJX9mGt
ITAPdymmY2djjNulP0BgnJZy2EWDgZUR16rZ5aklMlkgHHzbOn5l1KD2btClptpeHiMBcK/iImW6
bIu7hF3uO0sEK8bkkXsi7OKbjszaZPOpIaO+dMSqTcgyrGDF8nbDEdu619aMvTdQUQzLtqPU0eA3
GkrAqor8ReMp0is5hTcLFMkR5X2Le1QvFCxF54F8WRbdO6t8KUMEcie4owa73NHY3BOuS9xVY8nE
2xMXNTJjZmMA6Q2d7H/0wzjx3dgO0mA0B1kUURDbUPrrSeQMeMSXFpN7FaOogE3YekjNPAOfzneQ
umzaUvtOc+blVxF3T750ffuTW69TQDY1ijDMsD8ZuabqRI1isl6wO4Ddr+mDupOktNorVI1qd+Zz
ACDonSxfzqAyDs1CFElRV/++wHp87aMHwEmE85HM2kyBmd4bly6U9mpfpCXMmsaogxafJ31F3Nv7
uY1QtjnLiHZuZR8qlpyN44Q+8fcfFZiQ44Tuo2FWh494MrimOwP9B0FUMbL61acMuTHwy1Ek08sn
+cwCxDLQKnchpTDeM5o3h/UeFyu7as+jrP6cdmrkUWTG2jhxUdr94Kd83AlJjnamgszMvbhfQ/yr
C4USdmDPrDFM+YUW/SLSQvp66XRn6iwoeS2MhtJZ50D/iMFGxnVoBeJ3UXs1urAvGNynH1wQDLlh
doX7ZJ0ld4oJHBp6lU0SzOIf8iX+Gzc2WB39ehuazgGiACSlfmus2AqqStr9+6InGPiBYdJNM2Iu
0SPafA5zZVd4Kpsx7iNlnlTMEo7I+OvWIga8oj0FClcX9JShbGY9AVGVyi8rSPod2qllOhdv7PJZ
WCSkJ0fpWv3jiSif9dVM3T6PXWIBkc3IALs4UpgW7Ldqvdf2Kk3zH9j4gtfrgm9BCwYCbGxvDV/g
xcEVnTHF8VldrOqRJruQMu0vo2EWZG7nCju10seD+Kxp2pbK74FZpUbHyWeW1YxspnEydFxeCPVE
SK1bXC7ron67oRVbUL23kbOx1DEhmjEdsm0D4P1xBDVOY5UYA9FzX4Aec24mmUpS1Sxea/TIiNNC
PEVbF1AmAB4XXLCi1EP4UcAwne2xge06uIbtxaAwwBFvILGO8B09nqDvre8hsVfBuOdNOh4tE3Tx
mFn/C/3byIJBSAfRX0rNA1aawPmLsPmkXX0OWX/vo4XEdt3HXTinba2kjhTK68pGy+UMUtcjy2AO
4cPthkUkdvLh7Ou8a9MfVHR+pTDLQRnCMHDPFMjLAWlkAEsKCxKW1H3y5x834xztzrITedzVeqjU
X0jK+jBFq59zCUP0NwOBQdpj8XzH9Ran32X9+4OBvoG9kwoC3mMbpb4uMYN4OMYEpB4EK+GbwhvB
Pe0p64YwKQ+A7zFApUY4Rek5VeEHXq3mSelTtWL/8nEZrp4oDMXKJbgVnN0Lg7hXrxPAhQTOhAGv
OBhHiUE+s0kewfLQ6wRVeHtNwd0dMoWJEAxuyk5H5tM9khbNOE7Fs0YB9TTWNrJFUBU6k7qf7C5T
gow3ArUmyfXRwJc14pj92L4HnPsQvv5f++uK9sqE6ixrbGOGN29McTiwnv3hoMwHiI1A+9vdeZOJ
58725zR52PGTz5VdZf7Xn+t1gkPHCrQUjm8pUx7/OGiPvEUyIAcjt+r+JWpv+ot+IemfVHmGTQv0
USI4px3D0ZtwC3DBYGEQ3EXtUIKIM59tOPIYAWxO3d4Yh6zOXn+Ia2I1/cG+aTqdwKdE91grqirj
Bn5rlBwGFuuOsi+Jg49plE8pH8vwIqVsJ0yK0CwFIcOukrEYFsiw6SnNh+DJ33PHIoNTjpetnVK/
NWVf+d04tdv5ezPv/oeo7GcZqYv8dcAAkqDtsg5n36FPsYggsDORTbjqJha5P+8UhKhEphwonGY7
25pcmx31gX5rHAIf4mwu+X3iohZxOYStenAR1e5DJaEXgsepWak/pY1YQ3TZ8Bj7EEX784stqLXf
ufenNNT3FQQhZa7RQt5WvaD+QJqQ4OYLb+sc3jqiEBU68emW8ewTZ2atniQit51+nhMyw3CuXXDz
a2WvDJD1wywO3Oe8baI6UvSXjSJKIq3O5VRfjOvauZvagwRYOEg4/xBVukVDWliOaxdoR6SN6y7w
IIJzbtWQAF/YKEringJHfhtwCuT18jA+khtEf2UxZ0s8lwrGe5vMB4eH+z96MSMsHBnzbRGZ0dOO
IlZhax/XTuxSwNSb3LL03B3/Yjf9Xfp9QfP4nAnPIdWGfabG+EW4E7Lx2GsG7o+LwGIUurq9YnCs
E4jElxkuTZ9uuE+kJVrm5YAGQXanPdwu6Js2EYNrH6C5nSa70q8PD49um9mSgAbPBVHnbjRln9j0
gYYaStbC5k3DUG5heO4y5DP49SH6CJoGIHJmlE5H7hQyvwPeL4+rpXgGc033/qnmj3lBtk0BL/Rd
7bgtCQASMsr6B9wnMyR+JdFv0YDW5faojxGTnqow/XTkuyR4ERMFIigxxlMACyEt6iVFdfbX3yz9
TvqVPhKoS/OQBzrZnnv/gSP5dEAPHkL2PPlwpHxr3rZUVciMSNsl7+v0mKjQIKhYnP+Gn++CR1eL
HAnrHsLA6NLfE9cPLmIhUsKHhjtjluGMgDppdz3uxPZurrlTs7gFK5li4wMthxOXkf/7Y0E0DeP5
EXTOq5nVpFal/1aEFbJAOTj6v956EG1xfiaEHPi5cnbtzyqpUOVWLgOYgeGkFl/1mj5iHQUHbnSp
CD0Z3FoiAHqR8pw/D3fV8x3rQHTNR2RFSZEGeE5d57ZlRD+ZNGMhwCykdZGSs13eZASNrQrvXl58
mGNIDRMTdGKADcfBxtK0K/owhzWeE2T7PNKktZihTwf2YIGUz9jgRAaXFf4cEJoVQJaDfZDkoILt
tdNnFTE2pGnUp8wsJLMWvw7zFUWTMqN4RThgSGbzu+BAhOqVwy7kvF4nih6PaSsjSWb+kCdI4ySJ
8+xJ7a3keaYb1dhuC9uWIk0t7ZPefyzRrY+I5/eeRK9vvk67Z4iDnBnhwrElbIhB7hKlZnr1nNVS
j/DyXlfSoFfIUU6IPCGGqaX1PLdCeG3/S2YMXe/4AM8OsYvk6FJzXB/w/nCtPeJ4qL6izsXTTDUq
W29NhREMBFTjG9ScISKjV8SarxkUonul/YAB442XhpyhlX71qngFXdTnRlgLR4wHxrJAdg3m3Y2Z
Cu+MNlm791Kd8EwocDyD3OV8wunOPNlYJQKIgEKvLGaqTOQ7os8J6bJfq9PIt35HYLRKCj2RrTcX
jiioHqAm6bxwQbEeHELoUVkx0sVU0Vw39Sz/SAbJIejcQHwY5qwE6NAgMf8qn3wkP/BS1WV6sAy9
Qmjg2uGCAbiSHPIo7RTdKKwYN/qg0oEM11Fg19HWBl4K0tmamT6IkXhJKM9RW+ynd1kRFrOhN0WG
dWa5zSna32YgkeqgRvE4MQoA5o8K5CVMM/hEHM8hFcaKFRSPCKESwMF8aopSCQEzxkbCHOYLpZHx
C27K+BKhDHo/UK3JmPhBTIa5GEtIv+2YpzPK/z5fbWOPOkFdM8c0KAEcsOuRQzzmroU/GFE7JF7n
oZDf2BVNSKuDqqImY8TAoeOZaeGswQMT0I8uc24YqkAAY59wKbJI0CtBUAn4VDxNlOzpNlYH3187
6n2JaIgDEIDJwvZKf7sRTt4h0q2lqgzybtp4hnd+Rp1MDRQh3jSb5rnbKG4nrZa+sjgMRXjLFaVf
XR8850k3L1mq/qQMHL7bbyi6CyIBnRY73melOq69RbNOhgsYhqhb0NVd4YNYzAN4SzoU0GdG4w7O
w67YJj2Yu/HH3D+Rpx7V0SBngUFDod9dnsR0XX5e0jrhOyJejQYnqUh56SnwtSpzOgAOtu48nygT
XKSzqLe+zU9UwnHkH7hqaQ7NoqFkHn1q+UHXbEFZvqpdFkEKKlN4PloojD4o/gy6TWQye9g8p5tY
mht34ztRR6JlgWR0hia3KFGyqilz12/trR4d8wuH7X5EhOdqgxI1KXC7+wYOfTZFcXjy5v4YAupb
kVwcQ8a6geHDedTVSh/fH5y7cIjGGtfwYNRTtHVA2Y3g6pF96E/a166hipmyBPHYmE8BjC701u8W
7hjWuCb4VkiTj6oArQJNDLsnGHtlP0XHFMmhdEsNQEUlDvvoZE6Qz2/1SKyfavB/4DVtoTQql/fS
6E1qu67nV14Cw+WOjA49iMVPJHCsLZXSDb4JlIICpxgNc61zzggzGIHGcU0emdOe8opnn+xfH5ar
pVSZTLs+bOb1bohvI+9INo5jVuRahGOlo3I/NU+KQxSgPM0LBJG3Eir0nyil8Gr34qLfcTaLiB4A
Swe1EULoEgDG0jid/w5blOsZb+iK89piTdZ+uKevGyER9wK41XOPGGzdn7XwZ8V5SuxcCc2OZ2Yt
TKLVisbhquNI8gH4OIUQw4/FLS72jQsGoDCFGHk5LsgzWsnacXaSxuS+oIVEebREn5WCX67AcRht
TvcGh4lh5DvxRzbtog0X4LOS/IFp2PEJEsplOCpkjxc65rvQdwdF4PyYv83lZDtrwMrgNShMN+Ix
DyvnNi0Eig+yGQi6ZpxXHn27TVqwhLcwnY76bHLwUe6fSqvX9n/ZZetJo07xUAtjEFH9WHern3qz
j25Nc4W6QgljkQ/SGMPZ9fIhMtVE2yYI2JjYACVxAB6n8zck/Fu+nQVyz9NMqCo52luy6A3vSQuE
EYimZD0K8JoJu9q5+mKW1y3LZLaTmO20osJ/iaRQllXzTL8eMtfmuCNs7OQaXaCm/pf0TTS2XsES
6eXHhTGqFHPLwH6RbgKYkpuIufusEfCw6ZLZWkiFLtr5jhafnqOacaR4da8gpd67ymzj+u7FYovE
TA5dmGrMhusJcNJTYm3l6LVtuiJMtg44N2sQTj0TpZTAcweg1mJYevnb/vH3AW87zZ3J9/7UFK8G
39ca050rHDnXriK1KJwn+HnMPcdCGnOrm2mBk+0piJfAdJuJGWxodBYPTUJwuv/cpDHtVUH5DYSa
NiwdmNJJgKNJdXR+vbb7/zZtqO7mMa6fDzhy5Xn9enTI2mO8MAqdHUrAVYQDmnyUOrG+nBecpvhu
ORGLY1Ed2BR3/1dMJ59LZ62WWYA7fYN+RzcMbt1K7q249x5vRFo5CK6uMCImrQzA7+7yp4KPFWNK
QoOlcG8ep2rQU5unN0aJScfBM6u7qO25dIVM4k3Yi+GcLgHjLXKIi74w2N7wIRtRze2sAROAoqB+
rnlra+CiVNqwdLQMqPWw1qqbqsk1oZU7pc6LVehHIyTf2SsSmILEBvsBaCb+B0JWvx4EgeoTWQ/S
aB6qHIRm4pdWBvHAquKZgPx979EJANz7p0Wp8CTUdiLHIDc/ZTfMKV6YXQ7L3ox1s50UNSiNt/JJ
4nD/C/NQe5r2mf+MXL3JoGY6LvqOLJMfh5rxNWO0XF/nMZL8kNa/dGVIXu3Bq+98KdKmC5rKL02z
gwYamHqQ3TR5LVfyapgsXrKsKdJmA5TEj176BCaw+AkFawGpnISjNj6wjgFezy7OqFwpt32hr9fq
Ap5lu9kyBvQlZPesQ+5suH1astd7nuKuwMqJrKRcZVawJftHt4aIPBGY0JtNiOqR6LJvlwuIt23x
WdG5hBXezqQTP1bISn/tKQgWwS8VxHOhud0yYKaxnzCoF8WsMCFKN2cwjSGrrwKULKXkGQe3NW/l
uRmTLhaRibwTsjSTUjJMSNfDfYX1wdCgXcQ3gmFjVS95N22PFOHyy1w9FUv+TBBr1mlBwzYRTuGK
+4loAz9CMP0mqAsznZ7lFgC41wj7PlxNz6b/Yq6DKKlzH8+DL8qAhLcRm2+u5l3McOlVJFoOqThW
bqB9QKOVuAfiLdpNN7CUV81Sn5D5k3ITaCMR5SY1caxQmTDIapnphlf0JThXtGnlXpWkKambVWks
Msr17bJDKZ53ogTeD57VnprD4R/RLakwRNeigE+0v6dD1/XL+vsDOkVpwYiNJY9gh9dyOKB1nuoX
VDPBlHVsBoModDoCRZLRa8CpO0aVe4fjFcOkSj2o86CHdNTauS7FL+EbP0cjUmHumG2qegnAEEZa
zYAme/8CFFT6hLP7BVyPzUcffNrUv+WN5AyoQtQrKA+vgPKkp5XBW81V2Wfn+4XEfUyFC5za9teL
OwKlYhjB7fKe6laaR55pLJRcyyvaSH83rUNvQAYiZJgnZcNdZCnbpiKZsZjNbFn3E+VvejOXNM/Y
foPHoKj028YHgY7i8hV3cwb02LKGiE1KYpTiLOuNnEClTprRlmw5i3bijcwNqRUJHaPEmQtFTyGm
dXRxTw1EKx5vLNSREX2DCi3y+qf/l6n9SU2PCzHId9f35gkbFB7HoUkSLdEaly5s/5Sk2vbwBedO
CY38z4wIOkbcFRAyyjdXUiU4/SkbpVKCuJdOYhDV3jO9L37ry/nPez6zg00ifvCiW0hnOkRDl85m
HKZlkwmqZidGx4MY40a84svzvjLOw6IdNHSibf6ux5wYlrwwGRfSywv7IwN3spdCL4EvqFMOjiBv
lR5jZw8anRTjKaH6ueH+Zv2QZOQ4xqKpomP5Ma3HZWCovi1iKtjVnxQyPs8tMqXlnxCLafcw6l0S
jxZlxp7PtnrS0OX9BIcui+vRtqmjDLotkwHiRKbB2DWxDeQjE2o6q1ZcOq393hZbtSE5IZPHd/rU
L0Rmb+QAolkRWRvhM0rzwZJxcZB7iGdMjwRBvwihVAyYFtil0zcrWSnzOSnAoKPk4o5oHyCDkV/T
cy/vDT6vp11Z/7e5uNR+XWAjbphF5+WuX1pKtiljewX8AI1Yo1uhrCe11Z+pJOWBBBZoS2MZWyoZ
/RoNtOug1dWY/KDN/xr98P3nWnhkLKFkSNgE/DlXcZMLC2nEHzWS6Hlj9Xmp3o0rJ9wCLaLrBatE
49OfRIbLlh+zqMes4nDMlhdISATd5lWf5YiWfLqKrMDNlppr2BzXCwmXv2JWmAj5i/UACSw8HjgO
mVFgdPumzokI2G/9DjeYneDg6pvfM5c9roELyaPu/RlIcYgXSjaoeto4N75tew77MjIEJsY1OnOa
d6QwsQSXzdU9EK/hWly9aFadpVzxmQFDgJkB+bjiaKwOivtfUF3T5HrlbuOrXVAPIOfh9Rm3NQkW
IwlGoQiamKsgm/zr52vSWiOIW1nmemhI1FqNDEaGBnaOxm89s1xSUT2fzGMF6b/9BsAlLkeWEtnl
hZSzSUJUvVAHUAQO1jjktoVUBsrvVC6lB+ABA3+t/fYiSFkzLiW/nTuejYHgGchhAEM5S1HNYn9q
swmffTp+s0jF+afedtGQFn9wrP+WR5HrRxb91+7B+Izv1L6mIf/eJI/gqBoPkM6ggfr4XyxYmgAU
zoaUtG0w4KXXBgWhvYD9CiXJpkbqYa9F/baKuP+InX0Va7t7bBvUjzP9wkbpCCcA643bhnlbR8k7
NNnftRsP3jXp8OFqXqYP3XYtVvWclZwOywPOK3nOefD9L6s98KjOQl3cSai2yPeKtCLp82c64shp
0WkSomOxbnjWZziTICPyBKGvcdsZn+uYEggt3vLXatWG48S+SxKVHuJHe7bBU1tkdNyRHO8iNeFV
5WrfYxnUmHTlciVmg3S7Bv+THxUXmo4t11t63vWEZ5ZPCeV6qQWVo59MfpbuqdCmi3DjUCv/klwS
Lchb9XmmIoMjn+Rb5Mk1CWsF7G+fhE+E1SDnUzSGzAdVJ7PqRvDE3aN1hTO+i8VqnU/JzgnI2PfP
Xe98iGwUm80M2cjmk1v4bcHe2ReFBiz1u6fz7CZnBYUpTN5DDTehpuWatxbWrJ1WPtDLgTtkc/lN
aUwUnNMiqoReawameYMTKdJzda6aOqpxDjpf0P32ezTix37EMqLUTtv/iQ7kjLPHDXDPHVovLeEk
LK/NPq9NxVBmBjchinFanxsrYxhPXPS1OsUx8pB286JCJq78GCq9nhnydUsDaEOWHhmGrFBAo4y6
TxvK0rM78wBRJ3WnKHfGdgLBWM3nWomSWdiEgQw/RcS4VY4BVE6kPavN5z8efsEBVVWCIwJVw1po
pQCO8+JJWD63sDYzgDc0UKay6M9hhfuDhVm7FmG/SvieaiDdUKvlh+TopCux/9UOoMJHQS9oUK98
YYE6pSw54B1KffwKf63ImSiLCDYZqPZ4XgoUY4u5MvwHZ7nY+Jdoitxi1Ns+3xhjuMVXOJJW3KzU
T+9jt8j3lHV4gwTELUj0oL0Qqqh8FeVY05iPjLunI+bPtsFF6E56xk//xJ5j97sWrotoB48TMm43
CmZtZ0OVEV7UvHc5qI3q+XZ0FVc4nHmhJMCGbE8tGwG11Sf7sxf34UHjvU93zB+CiIni48gHWu1k
5YoflM1YjS7DWu+u+NFf893t298CxJWdcUq/LDDuAlB5eXAVy/DPZKUDw3KGXOib2ydyareOFX7v
uQxgm6wvMWXrbfYmCXekx1WAV2Nty7wokA1f1DuWBpclpAwmKkIbgtb3Mxhra/2TpktvVpvSHrYb
2WgJj7faa0PNymg7/307rXWgh9LnBOYX0UUqtjqBB0sX5F40S7p/oFuuj5CGWNULfDXTHs+UNIzN
K8Wl1CyC4DmuY236/UX1W0Ox0LsYE0I54BXl4jYKQnf7knhR6ffs/YGum1C0K7sJzEYZX9XzO0nd
vQnphKmxJkt4ZbuLYcwxYXRlQeVKfFv2+RNgSOovgAsRtXVskJ2RblMmQipZF4p6vcQ+SriMaAHP
1Kms5XZpiJj4UhSoCZ4qwwufYVM1s1frX7aa/FiOqfyOQlRF7sCujTHSPI/oE0/f6B2k82WuyNDB
LuUYD+M1Vei4B3/PDt9x4vaA3pJx9JlV3vNTAh19EJPHjXWVqzLFFZnmSVlUSAG6CVs08OapFOdp
oCZwL/9ixLLxf2Nhi3RGDglEiULb+rYgTWQFroQQBgVucyIFBAihE78sTtxyqwKZnOyD0bwVUWSt
ybILiZiwvOTPtqFwZLTg9BwRXUhShdzfJZJ5sA8WRujPB0WCQvamEFQdYa39snSgEuiB3JHpkreY
ZtYGzkASl712svrj8rr6brJclwUNS2hVJmiqtjMqoUScVff5r27KwCZjF2eJaSkdK9K2otcAP2D0
l7J2dbBp3E3UBV2g3wSaEGMTC17aaqU8B64fkwjhyZkI9KRSiD3lIPQkeZS8oQSVt6Vxlg3vEEVg
zMqPWDanPSCehXOlcukCnweQszYDwC1mO3dqlJf0sX9mrv/7Abkyq9CT53LXFxjeoFu0ZLHApI+O
walVu8ibjneq6UsyGu480gQlyQleLXi2oqSgCjWXQP/HoVU7k7khabEbZ/8oejaqu/VY2izkiWVI
yfCuCehToTL2EQ8AWnFjGdL/17vwTcc4kBBwUcM9RHZdUGXZLLqPHkvfbNQzNRbaggkzIJKjeITv
8fhCDdKGvlbfyvlzkbyubZ867y5UYo/ArrlPzq1oUfsCQL+SxBjyPo5+jkyIcOqx5SG2zgyhoEht
5L++ntKioPQsSZ8x0D8dG22KYmz7pmLLPZXNPnB9z2f2mnkjjb84l6s9o5IuTaQ9XZYtWQ45VxrJ
mxFx5rz0dfliD6nGUwTMKUF0UhmP0ZDKlBD61ro4/bm+7SUaXeORS8R3HMsLPLVlXxTSDWqlO9Pp
0m5Y9aRhvmtqbt4OyiWS4rFC2g1WpbFmc9rI2PAdJTPRGrIZ3YfNUewUibu44jA+clEwMxizRNuW
uHqTcblnG30wt8uCdP6RwfDQa8vu4V0JV7gWgEzSyiWDGGK2u3VPtTgtSlhARNrHbFVoiuZ984+l
lK7NtCaNJPb6bfnLb05H2owQC5a4vZ4xf9NJdneMq7qjsdkPaBIinC4i29aIi8TJW+uU50HTlvoV
ao706qZKcpuQ9ED3mLZ02W42WK4AKAbhlvx2AYWDpTGOgz8b7Nj7qgRBtaKGvLxWOOZMFou4H2cj
3qss+wubK3cdIfa8DotRZDqhsi7Eg1S1G17I4driIcobh7uWkYOxzjQ9ntvdDFPvGGfCOZ/1wKv3
DMTIReLRCiaotPHxprJQjfOXcIbxhJDwT9RjiP0IfTkMQgpViMubpvQbMLwTutb09DMbSj4DNRqQ
CPwkBeMhCDI4JtZJaKvlw4Q5cR0bP2tHbkWrD+mo36IePtt28NykIsPwTlKDLIohQewSNb5ARFHG
QAm9d4e2hf2Cljwn4hD+nT2XPpqjcRnHMlakVAYINAsGO4Fx/IqPPnpcDOxdQdbVSGwg2r1gLYpb
2Z/KTtkHTA0xIjIqbBe0tr7fhz8Fh41VffWJsWNMzLKm1SGSqzZyHna+wVjpOugqoLRybN4zg5DR
tuScLkGvO+wxZkIFIZSpw2dOyNXbs5rZT9Uy+zA5x9A5GG8ttd0oW3kWAKV2HMsEt0Myp2x8M66F
VfxbdfHv2Q6iy8dyuR7qTAOXj53VP+ktAV1INzW1Vb02YYZhtVs7YFoSJB0WWFT4VK0GPTFAoDbS
h4PHOJtf8UJX6dTwI8H1mj76lkWY6PBWY8z7h2fM6mnIWrb3IP4jDn7Dvfkk1DT1ER+Fe55jfbLF
LT6rxFT5Phqa+DQv4T3CU3Eznq6RHGPisM02ktBSvNfB7bwMPNfk/SDldD7SegTa/LVvFrR6p056
quqbIzsV4WZ7Ocq29rvok7DLnG8TVPoQu5RfCASpJhEJD00QZRoRsWBDNx+nB6ngq6XpnbIIioD+
S36FgdCb1m/n8thqfybIbIX/UgrtLbBGUnZKtBzErwSGASuNd39eN35k91ddyXsrYOQXrqWBSMo7
WhtaaL9An20m7DwQ066StKb5hFhpbpyfiFdWdhYhJJ8Bsr1J2ZJvK8iIxkEyHm6D+3yFGOKkbyf3
EFT4Cp9KX1uXyjEGMNKCt7aGJ+ebSldx7zSecYy3sliLSnJockLjH2typbYuvrTevwLU7sj8rH7S
Vs7VEBX7txIxD5aJrK66e/0Xgs/nUhkho9Rkr4z2oFG228fwc/Z7rgPTRS7ucS8G+6bvllvOI16u
6jOt1X8ZsZKmAbGmJeh5ycX8cehIqCpro7f3I1LK7QZEST05NBC0tibK1vrKHka1NBeQlmOTWEUS
yT1/AwdCDkPab8vLFKZVFP7MGmwEDoJcfUDyFlZ20qwRczm59Y+1ha824z+1AU1q8hdHHEIkIFyq
+9dg+Gdb5BCpHY5bDCvy9Nf8OHX6OcAFL/Ntu3u5Uxu4O4xUASg0e5njUIgBxtnmvruBg4/EfEer
2NxFWi9q4PbBNpageSGpEVyFba/3Fqo8rjb0vp0nGD3lOEaZn529PebfejZBZu0b+ASMC1++h9oy
hiP47SvnU03fy0YejShMCfPW4bVD6Wg+IxDS5wRZnMcwT40dIFkSUudhCt5N4yMPUK5kG0YB9EcQ
7/E+o5yikynyUp75HwjtaYmWwuyfOMDSvX8sOsRjvIs1Ssi5a3owrhxynCgAIJztE2lEgQnRlxxk
HwskNU5Mh30vd8s2dR2P9hqR11wtwBbWRWF/8/zmMJ8sj3dV3M6uye2Hi2L9DO7t+oFizlgGBnle
sVNgKvJsEWY/g6IyJ7ZA4AB7XDwbkpgG3AG8WxWPhkkKuI57H76Kxnw6nAqoi6zqxOJDjp7LQ2Ng
tODMjELlnJbco58dBkTDIXQ4MmawfaVWlw9LUyiFVE3bzgYVg8D8xE3xN8VD4x/Ba1cbC5RL7h8U
JU9zVZSawSUmz/azwLZtPoPwwBB0gMObKQiSk5hJ+YnC8QI26ppwC3pLFmPm0/0hCpM+NoLIIDOm
WNTSII0+C4yAGUraKPVc9bthvgXrAnY6eN6o/8yNKnNM2gWjvWirQHijgiOvpXY3j8cC63S6ureW
vUsCw6J/8KEeJzBokRjlAbr4Aa32u9EbDb0lJOYb6Xb0wlC4ysHdSqp2PBR4RBbprjRYtS1i8Zv7
o4/HlsXYJcf8PcRXJfW/yltmckPRlMyqDhdkXxSrT2gmt/WqtHEfbmb+zaJ/WRLTVwxKRlAgQd86
UkJ74HDvm34yAnmG/iryTFyn7c3GE7M/eLo6Nm6eBnTey3nBQXHK+mGrhWUC4VbfZ/iUtWgyDrmg
GIKsINfhi8JVsYW7/Znznh2E14GXzDY3vgqvWStU+nhBL2e1bAAiBmZ3l+6PzyIRizJEKTH8WwMb
BKEpl688QcD5VCujX44jhZ8anSYiD64O4RkrO2ft0Pvkrmj5pCnmo7o36VruXaqqvB41ttvrr+aK
zgm1uRaQ0nGiAcK+1qNqNeRfBFcHe8vUns/I5TyZNgOode0pyDxyE7pidickMV07HRAXYnbOjRmW
w15T/xQT6Pm+6m7B2rMtp1ICP2zcQC+e3KMVdlcaKUk+KKTMQgFFehJqu/cSKLH5AHSA1UqHwX6E
ZM0eyp26gcZ0xxOFWQpMWsgVbElmWuciT+hYhKBn7O+BS7Miq/xXetGeixR1DMKjXQX5+BbnSmJT
LtZYOq8iHCsdevtS8uQNvNd2llXNTcRayhC3DL+EirdpDEv3PDmiRaOmlhP2TJsZNRlZn7VCKdvN
YsfBo6b4quqovwfrrGL4UYq++R4HD9DuJOh0MVxqPYjYKGcLmaL96pknbxAuVTqc/eV1jTZozahA
25AkXIyGkHAXLCkakUCTFbTu4pEft9TOgu/qeJVPGr7HBC0mhLYt3yzBnxyULDkq66jaI6kr2ywf
yf9yXzFIhYeFK18u0E3o9umvrmaXdO6lZ8xFf5MI0qcvJ0DhWQuR6EWfBRTWwf3DlBWwF9rjEv5h
Cas8+gRc8FLkQztNvQ1TAGPZeFyydWlfs5dw4o2rLHEoOKL75ib7VAfo8LQiGgga4KWKW5yeGECA
Eir47JO4pi74zd3ub24Vj/M11RXG8CdqWEtKv+vjpujdWwKlPEDVauNI14Qnkq9JdMkJiDOzijWw
V2w9ilmw4CbdquqhJogEIRvOyf7dV+TV+OTJxxI+RFBDAiOVaXUvTk39KivzS3mPtmxhDTm6imxa
wOeEQd0aNO9IFVFuhofsGz4hVyQ/+Kv1q2+iQ3/nYjsQ7yISrP7PvP84yVfbgReeMZCumVIhtW6f
UpHQUE4KncwbmbZLRzLtdkhiKitL5rt8qUsSmRPII4GVVUS/KEOxtVy6u2kyXlc2SLtdS3el2q6G
OaA1PgT4flzjQjKrUs6EwXIpjLImmYAdR3TrfSp22GpMknDf3uAdLQa1sKu5TwSwEZFuiHfjXoVH
TsuE2Vh/HRFf1Fj3CsrDuABCMpg5LOr/BZmjI8gaVN35gXQVS/wku/MMxszG6FjlDMb9LUTVekdg
yRT2RNr4adAFCiOfX+5+vpUplzjEc8S/iFDWvpcbRUT+H8BEUUipa2wsCLZ1g/4O7zX6FNjr/+fd
IqOACHcC5mi61T4PyR49UdTjXxESQmrO4lyxUEJ3U+pdFg9aSUaEeX4mHFZrg1pw+0RH4+L3yRiD
RS8QiOFKTMkXP3g7FGJveug/gMoT8+JMhuirY9phRg2nkhdf+sOx3IbAJuzyTEdpXduoN8Pb4wCb
mD791vYuizoDBqjVBWVhdM2Gz9Zp1M7sVUj1kSAatBEN6lxoHVwBKo/SXCZOrpf6y8C+Qjxo6zf5
pnOGQ0jdAdn9nr1j4N316ZroeDQtyjqRJMMsfcTXWyPauS7ff1Fj3C/5iFT0Yd5IJwWjSEmkdj8z
+iN8fqeKGVCyqS/jkyw6x2d4RIZWsvxkQqK/clmNSx3lIHvj5wA8I3qs+EAEn7MkPm2yMh1m5HGd
aG1SB8yTuaNbq5IF75G0KGmQk8oTAgChae+EU3plB+5klxA611EjEv/IqHSr1LEB5tASEiD5rBOf
x79V5KhDUMk3RWjaW7UjZXJzODL3iQs0SkcjKJ4M40+G2VyLnrilI9YsBJDVAv5c/gClYPHd40+b
EaTRbCOvKC/ujcTVXKv5Fs2Ve/f6ifa/p8/enFIZ4O9sMIrnSGzYdRgF6mOLOvrkZNoHqiXPNnan
Jw7sXyFS5XYWuScOOuX6mOwNE5zfMBbsbLoetdbCfos10LYaxNdn5fjjttPnZtR2jxwk5XoXhYr7
zZt7N4xbt0dARbIYajhVxEv7zNFT910G6Idt2Atilqv5D+iQf2+vT2PYSsl4sE57mWUlkwwl1Wd/
KvjrUJGVzBK1xWlqPOSt7xJ+PArcfgOmEJUE/tkFeikxgEyNTzGNJRCYY6FJ6uUZrV6fPXDtRXhn
AipmJVfNM0jDNxxXgc0b76NRFaiJtNXFwKt2Y9vBUsLb7iCAUj5CH3QwKwBnmaYxBOMNUJbMQzVp
P8wSo8qXqBYC1YXCgaxH9xMIqNWKtdwRFv6ISa5wOUmgctAMUZ0DMCmkc046/SXFXrk33sOIm+bW
2ecKy/NMFlp8rt8LiNfX1TaNFvp7qgGT+ZTTJAAbjfBtfUOxhi2tws/a1/0kM/EmgAYx7es4+mc1
Az08PUZ9g9BAoRvf8Z/OBH4aBI/9n0e/j112s9z0sQTC9nJAH0a9uxcKNz+HIsrQVEYlxXN4N2z7
b1gQOd1O4U+ulT3DDGdXXWwp3Z09rC1go3Vl0HYKtLG3wblg3gJvkRSYu6u+NcsJgx1H9afPaBnj
p+52hXL4u71bFMK5V6o2YODl8Vi3jW0lm6dseOaa3Ns0v0rDfUzZ9FccVaSs+MdMBdSl1H9FABJf
/HaM7c5pC3UlyqJg1UiIYukF0Bj2OUYYRoVpW7SpA0zg+fTHuPqHxxngmtq90HRPXGc2k1V6e8uX
BGDIA2KYluaDkndx76IGzfhNYdPhPyocCGIWrQ4TxrsD96CqM7wJ8bF4PvR9rxkZOqq4LnrfV8oP
MLL+4z3LSyu3Lj9fOHoGUE82DDr0CBVN8tvmSL73DKVhp9rPPwqv6VYC/i4dBiKvWmgqvInGROWf
u+EYNZae8jUi6XipIcEByhGhLm0qsRlcxqIsI5fzXfFbgdUKvJJWj3hPMu71c8vOvWJ013fwuCQ9
Mo/6Mzhm/d6+NrcwrcGSJqi9ESGK6e5qj7G/pQNiNAr8XzMkctGzu9KIa483tUfpZuG8R98Svjwu
iw4y6ZhlCLZDBfPX0CLXjwP+4TQ8Khd10skbjGEMffHVQiKhKg1ixKzfK33CFNlUSsptzl2qFEG7
fwYwRTWRW5mEZ4nyQFURDde76BEB+ll/1pPajwlFRF/J006pVBuOFYAbRrBDOjuALSXzi8Wz3wmf
97hR34GWEKz5vBY7TfLXmYOPgyMloqqKY2VPKltJ8Q+GnXkmbmxwcuuyfR3kwPgWlXfHrHa6r+0W
7KMjsNpuFhQJy130znlVOygW+DGWtXInnF0it1T9jE2RDDbHaxm8TqDMxPdv22yxaxCkpiR9l2gh
iJmwKaP1E/TVKWBg5RyPV+U510uiQRDXqKnf9KRJ9W5JkFYz+oAoQN8pGVM8OGozqL6PSVPVOOUe
edyRjljKbSk2lMVRYx/Z30gSAxzZpcwoHakdQbaSqwRqNyHDtR+SMmeU3wRIKrSrnrRL2v/p2kjz
cDBchdi7FSmx0zxXCKFkpX1DoeMIqHjsE3xCcreROZVCOhSnYvE8dbrhMOmAOsLYaYsE8BPmzrpx
sC3QSU+KqChHciCGkJesUxtnD0nUqxz4fcrMLXx2IPwnQq1KbnK5q/usC2Fq6d6lVQe3lqzqoyBU
tt/Q+7jR4Va5P21fLgmIKLbBrs/i6b66ArZY52Qv/bhHe9Sx/Q9aEOxz4MRC52+rcykdIw/CPN4S
OgE7SBq/MCB/JknotqXfBRxYFFL56116maYfeqZTKA76Cj0LQrPJV+L5ZRZtqxXTO1RwevGOzidm
F44QXHJzhlEG2ULCKhQkeIL5BGzRIySc4nv93csLjflLH9EO/QBSjOqmudnCu5eUEwokSQ8zVsWL
pCewDEQhW0TJdY1UdV+Od+SXTsPJaChkxnNLyW8t497lSWRDU9B5HfqKDLrDWbBZcy/ovqb2kT8N
mbY2VI9AVMjiwah7Z17fE51Oyb1L5GwzhnDU6bRQ7UGRlyqXWXwM0GuhqPs1JR326FCcADssHnDC
3VOidkc7cRPM/lhZ/t7RRQYsLULUe8wF0Bbh1ltf5EiCuqeIAWjGBaHjVEy+fHK0e3LH6o5dsaEZ
wd7JqfSaKFyvJp/yhYB3mZEZu5gKyR66pyxFsdXe0Gae8ebTG4fgQMotLeLqrOym1s2QF1iMhsGI
BSFCVZZu0Z3oqKvW0H6a98zMxzvlbpcNFY35p3PFAo9IX5oq9sSz0YCrvDRXIimtsCERcFgkehQq
xrgxNaxFUpAD+5IijGHzZ62QxXBBhXZGe2yAdZowSnWpFsF4ywcgO20qlrQD501aC0wtVOuB9xRe
NQwxYLfEkwMZWKw4Rvzo0kXNOAtSgcgtMaSnElB9sTM3tqqbaStXkIzhM4qVISxKmuoz3nfGt5LR
s5xQ24ab1mjBt1uydhYyV5lo9zWudnfldVJWnE678k7Kqzhrj16qSzHqFCGb4k+55tK/hD4rzJu/
UWPOmkxRy4bNJ/SW7bhkPJGFuXjiQmMjEpKYsxYydjO8uiS+2dkecXxahJwQROfTJDkexgmgIw6E
vMRxHncEjS3A2d0BMFB+qAzYuT/FY/VoKvWhk1cSW8rl1XFbmAaGWDLfbYXfZAvBg/7D+fnhvR5I
U213B77nOJExQsnpgM1CcFTR4VMpn6DDluVpep/Cdv/8C51ljQkuh1E307bgpCzYs5gKgekNCB8S
sqKpgSidK/ikqys5pBhj6Orsdw+8ikAmJaqW6RBg/0YgErnd/b1o2ypX4fzXOFasL4J1shB0h6xR
vR7lmYdtm2TM8qKHBq/atRxNjWufSJ/2vc/YwqyEmPNSIa0Plcz3d5rPdzf9efMuacgiqjOFMFs5
PwDtDRMbVGBim9yFj+jritTRS3COb5PebRvOwrYLIWjwLHIw1tcByza6vRo2zQboYZo8sJ3St485
C0gRfslXZ16jUcEEvv/lkgcpoimc2muuNMTAi8Thzhawl/+5KPmj4NR61MhbddqrxzHjxD+/Qflb
JAfIk/qhDpVKpAD512yvNF3feVuxUdJpcUUjxc2D8bPMB3pbgkJgAYrvRmIFlOWn5tzZziD/hFXk
qTEZlsrNMAYaL8bTkvYdesCcxZ885rinfAgNtTcDSZ+4E+2U67vshGnzObV2sYuo/I2uR9fteZ35
eJKXOucJ5T6drK8waxHnO6FKY5gRIxphW3Nm2N6NohhP6u8y3kCuix+Q7cZcZu/GuW6rYk9HfOKX
/PoeiYcdUSGVeJ4qrHYr8GSQEW6eRYZJrFOEkbCQtNYeepNGKB76caKZ/remlShQ5GGl1iVTkAI3
PbIiDtKnbPgAehmUmdAMou5B+BhGT1mOLbfTWTZIXG7xVv7yxLa2kBKUvt86vk6ac9mrrZUrJ5ux
WhKerqHs63Hd5jtHtH4MZGNCcKvvl0It/WRxeYrlTtMbxP+Jmjij4gb63JgMXSH/SXwHNDGxnbO9
tSgPAfDZ0cASiaSSWvenyeQmNYpsFIcKP8OQWxzkJmqm4y8qHSpfQkcUmFsPPPVKqveZKImBJcYt
l2hiJanxu+6KuqDpvqDMx86jcd7v3KvPRGUsByZONX03+ZU+oU5UJFWEqq5ZIUatbsxCribIqEGC
4bylWTliZV0gxfGg9tHzQfkcG+er9J76cn3php/Ulm3t+aKZmrEdHEDugwHTA0jx2Fv48wbkgeSs
FXoZONpw4ioNwyi1ye4PbDPz4KwoCwybyHJp6tDip6e+lu5dma1Kj641bkyp56ExJ0X6XCbmhrPx
f2GDBSHzLTgcuelblzKoM/6ZUabK71+tIgXDhJq009SII9pfq/bzcH6NueCZFpSdX96YplaNCYAG
c+MfuAtXQb6+rO9Ak9IksXpHWINcO8O1b3B6PvRlHVKNXRrv9Ubb167R6UrepRXZnMk93nhWYAmP
puQXIA+A9oOtWeIZmzesWhGg1URLTQDqReR+RDHPYUSYCmLYfd5Z2huMFJWJHcpLrz9up1Kk2p5j
RZN0GndHlu3UASpbcA8OljdxbHcGMgFRcB+QU4T3VlmkVRDPRbrXxhO+l6GNtotWbznuR+3nghPp
oX/Mz5hI3yXvy4cReZg0+kJ5Q9VbhYg45DicO8HLDdvItYz4/V8uD8n4UZjZAyL9sneyvHYOJVhH
yy3cxiRBY9tvQUanK6tWrRa6Y/mbeBJqMOOqpfn9vJL0Pc2C1iV/D6U+bIr0xGBfgXDgqFevSthV
g7kf2h2/7jXolWoSemltZgVyY+rSwFlst2HJfKLczLzOCRcHM9xD4g7tDqaZF69HPg+hEwidYII8
JPLhgpVVGQz6Eo8rBFyObHN5/FqJdrTaH9X7ma1S5Tsba1WN2K7obTjRZ18cN1zgEvrf2DU4g9Yn
qxWvw3w7VjVGFHrdyJE3b0rub6hjdT7VgVV45EBdvDF81mdzhnA4bBmJ/+yDtfBpI4VD/Bbra7Gi
3x4wPkfP867SUrZLMIDPCxkKv8BoEAl4yE4b/QiD+296CnNyV+1MHFDaKueeeb0/wSUdQuwMuDE5
SEwcWoyLe++J9Xin83P23NAlr6U2pFCG+JTWvRoaioRfZLgwOCbaNfGxJ0hMzE17Cr3Ce/s3+/Z5
nqYTKsZ/s+OfI1szCQAq7ehPHKJFR5KNzGre9QoXqE8k+4uR42DaGUd3gmi1/kIwGcBnFkD6CXaS
QIPrjOA4t0jPQmQSTA89PxOXV76Po6YE/UDwfAaErt5R0kbkrD/eKoEvZqC3IGRkeFq/EG1X1XuC
O1e21axpGQI1mgnAUGx/QYD4tSL4398De2gptY2cFP8D0dJmvL97IeHrYGAwz8CBnXvEFnFq5HDw
Uj1qIEEhZNSeXDHHSmPFFobN6BKeki6+TUVETQgpvTnzytNc4SQupwkb7HbBXJHJnXNj2zIDuQ/5
A9Yf5eaRkV7Jzng5KioRJLujx+FEJJZitGD9IB2leCBCJMgwG+VL+QECJG5gHw8N59nM/4eDvrPT
cwvasIQWNwDXKMuHbnkLmSOYXUWlqU33yHqy0UVpr4RPt4iZevyvUK+mi9DQ0rp9YcuvRbcpWTkB
fKLCWCczNOtGkqVkAhLKRiTmu53mQ8pw7TEQfUcd8MepF3fXV0otg5qj7/JrA/D4iTpOXt/RvCTZ
GEf5JQmRo2ZA+8ZKnbYQnjVJPau6067Qx70+tnfPMgclN3Dw1GhzycNRxCkdLY7iwDCysGaMwq4c
gE6Llum536lUSbnjmeDjf0IdhAw9LR2ciqoCks2K7NYGyCwuVRdb9WuAqDB5XdG0QG3OO4yOQWnp
cX1/R7y46LjK5XQu5q61jBDIuZV3ALKMcIxb2MVEGrV5LJLxrs6dk5kkyD9sg2h4OPOqLPgrcqoU
Db7Mm/27UV/qPPohlkic/EU7wRn/O4tJ6tqZrTluw1HBK8dHw39Ju4irtRhXfCplUb281YUm0MwF
YupMguePBCnqMhbrtjTw+qntE+UgwNgyb6+LaEm/NJLN6U8gwabAoxfD8bMTQHdFODPxw7pwYsIB
PSTzQjTNeL+bh/aMP8TteM9lFY+JHyEdTUBLPYYyeDrvM4kB93eGIfStUxk4/pLQi7TWfMDaNSpM
GaTJ1TyEO4yegjHbRHiGlEEx6xItR05+PW7lLaPhqY3GSLQXrXysHgnZyH80m9nbkpi3VKwEeQ3b
GYcH97QkOpYZzwNwqgzji9efV19LQF+lnnSqeszT/DTuDtE7e1Yxph6dGRvDP5Sts+ljvqlGuaaX
0GUH7RmgWn1PQohTEJye9OK93FNtdp+wxTimYCt0KnXyUjPgSF5g+B8UCIuJtdCyfB2Vh7hNN+9q
280mznTQZgyZSkVughhM6ffQ0OeYK0kBsYMG1qB66Ufeq5YQsCNiSeNW8DGRCdEjdzzmds8fY41E
umVqLNjIlP/UxqAOJT+srZ9DstRY3F9SeEk4dVuR/JR85pCmIpmu4wWT6QfePtTktbgOtDJpbF8M
Es//+Td4ULNJ7aREG+SHFKFEbzyS425PeiXOx/ErC8c1bI1d6k8gbfdIYy1S2ybe5D9xUunn8jL4
wdlppJz6miG4UtEfMfJYRglpyAam2fAlQc4dVdHwc11WwDFkXOekIm0cTXr5tci91OE3SA83VjPV
6ucmnJh+IrSVD7WRphpS2muTZmfuDEvOYkifpDDCBr898oMxtDmk0OCA//tXXim64KgNdAib0UzE
99JBTiRL3i+D3RSIFURfzQA09DPDRJG5QkX2CotkFEFQiY4GqJhIGZ+aH5o9JOa7eodrdKUm0CTu
l2oVhxuFVzqjLI84QcSqGtaURhDWKaiTN/jNRAxsZBlytDUGQ9qhHq6kK0sYLBgSJDf0KlcQ2rYg
v2a3AI8Y5PSmD9htWXlOlxCa9idc5XJxDOyRWJpFpknlqA9Q66E/a08zQLUNeiy56K+htZsY2dtC
HjWBAeGLL82gdCLbuvinrGt46DifYQHAqLsr+GsstMhtVWZmHvyIAsP0hZXZqqdku+DvUpxkIwKj
XFqq+cC0I3D2QJDsCZbW7J8lbHIJ5h68k7wJB+7zDkylOElLXdZlFIi7IxTgPC3cAm4EpDj6oD65
bgO0U41l79QkYGxZsFKuaX2o/FCfEMA0Xyj7PTthu391gw3txRLsoQ3Q2f3WZm8Y7KEpQRWqCUjG
hTWJrSMBg9vYtg3/SjNXSJspVc+k4LZlpUJe+zgZTPMH9ru6vG67+e9qQNnZgjEV3VeL3zdGNOOA
rKIS+t2YHa8SI8FoLLzZ24egzuxYTgJhT6c/WXYiJE7+7toQgRFVWtKTQFiap4K4FA18kNOScJ5C
1syg6I5pGOPfvuCXYXIyb8SJ1Oz2G4yjn0E4IzOsm7TxXMVAQwXVSMWtUbrVy6CF7zkqm6N7KU10
JLRtPfIJ12SG67GxUEpjbAv8d/03BFISTsHbTb3vkIsvSs3XvFzDQCkzLlmY5zUXqsXOI8zGCfF4
tMnxtvqAK9NTemuvA2dc5wQ9Ld1DZ/QDw4ZKWDLk1/PmZa2Ws0DFcXTcxGq6RtvCNyCCjrflq7b3
kqRaqeKF9wlqfkbaQCTaszk9Dx6zChOBV6fnOrundtgeUy2Sr5bWq+2VXSwmNJCpuqQR/oa+cfER
1i1SMY+nIuTrWZqysf7BuUs2t4los9WDr90x4241bHdCYKA44ZIel81S9I0fYVfCLBVCiSSJBOcM
7hxw7YQRoodrDosLvTM+fFMfuAxbHJg6hqansJBPkymQ9PUg9Jzohckl3tIxcLtz+89dd0HoT7t2
jWeuW22sH3h+82AwG26V5aZ7NVN1Et9BCMO6cDz/KJQNw/1BxzP8tA+D3c0DVANLcDi3svSqrtOf
Y5OpAXCBGjMAeV2Zg4azAFI/rORr+I7EZ/PcpnuIvPwX+CqJwCbXgS/i/UKFzH0ogASVGGb3RQzd
rJI8TlJnmGqjs99w/6p2DT69wTWKE9xu+yK7XBUuc70nZpjBZwvHC10Jjc4ldimihCEDLPi7i7Pa
BqFkjZxyGqyEWHfh7vUrmifZnN+SH3jaaY3jvOUDkWIgD0XIr48GbslgLhIx+w9hCtQFYv3D8zKB
2kSfib47D1xIfXJzFcz0E17nCLUFTwNnWMya50psW6cHUSZNOhe8A5Iy9HFAsZSOeyBxaKfMI23+
6YZW4PkeT572HRHD8CrhaAehSJ39haE7BlPSwYmQGy9ZC8z7uFjyqtnDs4E66AYZGPlKtVYHEAk0
zpAa75xTszf3/YWpvakzXw2oL0m4YTb0qgtwcqh8XFkjMrWP+UQVjD2z7wOqrwZxN0kX1pg7RHeA
3nqbirHm2BLl7ofOu/KrMCLfXy942vdOyHKiEZ4JhP+V+WRKvzL96tQi5UQLUjSMotDhWgKdjm4H
9/GDDF8DlhKxMnVDCNiJY1tvgd1gBZNIYWUkorZlebblcYRizzvh0lDnJN3kMxXGur5f6tERJ+v9
ki62cCEV/8k4O6aE6DoIclPoBqu5puO9x9ID30UrooyWgOQUnSLyFA3olfweKbMIPCZcCOSrhE9K
HzsHBFowNU0bK9lRgzdKx+dQlLQZQ/BGEK/tInw+TvESecZef/t/UTwZRKne5vcam5iTqdjlOxyN
u1lavrR0fWClrbiLOv0PyxzoQzVls1015AiEzEjTqWQd06BzOUis3ndEe7OMDQkjrJ2nk3HtUaNx
rz5wAbPwd15KeDm7tQUvWLB7DfxLoh1xPaoFz74lGTrPTlikQZ8khiYuT/hvSsu5gZatVFnofT6N
Q5E9vueEOR5v1qtlnDWX4DS91/jUABPZAbV12oa79zSRN1SBF3S8R/IXT0vaep7Okn80HEe7S+F9
Nekm+yTdcI7mT7RpYftqfQf5dlK3gDQHcFVLdMag2R0kDGasLEGxaV4FvxUioZjFkXj/Xl3evJMi
G70Z7+4F9mt6Aq8nIKi2O0QJ2f2++xIjUWqreR/qXfUrD73wd9o2iVVSdkMno5MW6LkUn4gBgYRY
CZveO397qLER8TrXR83vH6XP8AKnLFA8dklyD9J9D6u11nAVLOYgk6rQKgoYvyfEEquNXrgdH7WQ
/sYhg0G4ZpYj3DzSAb8+BO1ikKtMO/2+JII+gJvpas4sAoPv5xjRhfMKWrcJzj89USItcmc9sBft
f0Ugd7lvLXbhnIdQiZPLormjbno8BXhg3B6JIteqg3CSbgrLI9esUwT4e8b3pcEA1Dqt2fhSNHUS
QSTg+Xd02IsLkBaHfvoD+EaS43giyMZIjeD8Gw/zAWLECcLQfUNiQeaPGVOFNkpJ8r9/amSigBPL
kzCpJlNIa1uaQ8B3ysdxxqYZpPYLLz1ufaJ3VBTk0FZvpNNVWf9T0LKPTB7ktCnK6svnRfVPoDaC
l/IJUuNq/0aMuLh0WLI0JSI3PJ3mgjugtAUKDdQUvOSBNOU3G3/TzpBMorJ4XlqoSgW4rod/Oiuo
HtYojNctSfQtrMs69kZP+Hgj53ZgHY8emhk30QINWUSuI8JhulZjfzi8jnAU0O+KcDrPj9Z4jadh
4hAYooL0rkVuBI6s1+IKVwMgSnCo/XRqzYVHCRXVMuw75/L/nbtmGl9INR9UpjcU/+KbN+5TrKXD
sfo8sHyqZgUNwgvQSObIofb/ZlkEdH5xIuwMQ8zw5DLtY5MYmgZkq30ThpBv0a65o0AKHSukAnH1
p7pr/jqWNc267l2410BEYn4zxbDMsjNl4k+oRw8qrzAPuGJUh+32r1F0aGhOSrrTeHasK5dDkrYD
yWJMjZl+5moCxZ75m/hzfxDHmJlbVe/byC2jQJHn576qpTf+I7GJD2iq5QNFt+WPkcpBrvBnMMLY
G6Ea3Tcilgc0LlwtnmzVYzYLEc73w+bYtbeBfcnttjucbl2wta42IWq1k9w9bMtz8aPveFqvQhvP
VdnbjLw6wPlULfI8HuJs9Er02Q1mbT4/lz53xwBMnxkY7Wid232bP8N9WlMztjvW7m4d5WFtY3/y
WkzLF7Gy97rx0XBCqvVMfRyqUKgDuKKMClrYqCOA0I6T38GTMkSOgJP5j8vrxiQCXlBJoaNLS0sW
2tzJTBvr9w97K5fuH6/9xD0FLcd6jJaJF7kP3xVLIOV7MVdl9LHGtnWInJg/M7z5pfdPyj2Yn3P3
ijKRFFONvF7cuyD8clLysnPbP6TnysTXQw8IrOx9VC7vNGMmLoCGP6l3uJsqlqSwRfOpA/ziLARg
jE2f3H+5JPZYPCT/F3BtWbGWdMm6OBCAaSZa3RrjJPBHcKsEHKRGEOfymXMGVtNnO691BPuK10yT
PLegcnGkHXEiyGGSma/Xy6ElpKdZxNWWKeW2jDj9y6aDpJdMEfXsdmcbXJ5dmFSg6UI4FEUeI47M
VXbXZdJqW690DeHkZtMv3mHygqqoVmvq0YxsUv6f0M1TYuBbf807pIpH36DGs/kYyV0gTePZXQUB
V1HS2KFdFlusUcEP4tcQE6fPRLt6RX/p65lvlhMkG3xugnx2L6fXUGfyz8RUCS73uj743HSfb5Tb
TVblD8aeJeQMBpu4iBPVhEkmtyRCVwRbluFSQLbKNoo7M1m17C/FuJnHBPrFVhbiEjDcYAgkP6SK
Mn+Lu7nkNaNj+a8ioLD8G20Mhl6SIjyukahEDhFYgj+xiXS/IV8+Lwgu2wtK4mp1IJr3BihcoB21
IzhGvSGMuMdDughGpdJEEc152c4cJrw4pQfqoJHGdFpaeDZc4rk8gkRI23U3itJf0FPbTItXblfB
oS3UqfTqz0yfhbN2gxMy+6VAf/TO7Ho37EYVZ4AH9nOftNmvgRFEIud8i8vgrEAYsKvCOuPfAJy2
5QhVFKFIIH4pgs8aegxcOMr3ePQDk2j608SMYKYUmbuNOyBLosYZ1HIZ1v2bu5772CKDO9EF5xf+
Uo7nBK6f2CyihPqAfmQO4N1IMbhkr44Zwo/a637p017jT/9H2T0jB/E3HkrfZl8kcl0W8JEdNdFB
zJ0a/Q/quaW7YnQ2/Q9ylxtjhHD4sY3DGu4ITRW+oBzc39nLEClnzqmOr4xwN2AjxvwtcUh33HKh
Dd5xtAp2MSmXrptcI2pUwXdXq8igca/cK/F6G1+SCLKa4fvZk/ng2ZK0llKb2uivcqVXYoSd2IUO
3NJ5koJ6sjwrUYT7j87Gloyot6+JjXMnEGiGg/fFrd7QKvzyS3E1OwYs69BpxRzBMb6yRwywYX6e
xq4GynKMccuMT+NQ25OfIzef4VH6jPGKslgMkTnbLb8QzEgkR9cbNTdhWQyqcAbrr99ZUPnVAAPX
jgALm/xyfKhWs6GqC9j6x5mCard0RRqaeC4oioGyYWAkNRqnwWufVTPDKjnwew02604m7yJGSRIW
9lywmQE2qOtZay2Gk4jh0qamqGZYqrf52D47XL32suj52MpeDWi1U1J/Hp6HdPk0b9nD9idihbY4
XucMla/YTPxtSq/y2GHe3yxru6m+dnO2YLrTuCeGfEj8V3Hm156icKdOV3fDub9PSggsk/F/GV1H
UE07CuWM7S6zIbI6PUMq4bSiCNwwUmgnhJReK1dxg9xoa4qi+kAyO44/qVmGG6Sg0hWc+A7Z3x3a
IuzhFwqUHcd6k1tfh0yeFe8NLoYNOki9fF6xoVmfunnayOiQ3sf7weu/ahnIrDW+ONHuqed2MiaR
7gQxCggvoFj94Fe8TSBqRWcUxuDgZbSNNXzmn8dnbHBqSJwf4g8PdOrKWaQqTVlHog3vgbNlC1lG
EnsqCuIEvEesKmntWHqaLnXWo5BtVrgvQXFNwfrQNz5ujRCeVtYH2hySMS4Drb3Bl2sdqCUzRk6x
9nhcvvHoMGxS0Leuw9zyw9BxcP5zMKl9zpnKn14h9YSxWZRldc/tUhkakNISnH93LhhtRFt5qJe7
WPTT35zNDSqNWKiD70I+PV09rNQ9ccixLqJcAxhZEJE/s8+xPB64SjgxR1PBqNSVUvuTVJ9ph7Xv
E+ANWxgjITE/QXNvlyrui5fwzH1lPGmaGlE/at62oXLgArWMCoh8iGpl0X9VHDSN6TqF8RH0GIY+
k1EMzX6SzkvkEz0TJQ3+CrUn7KKayIpyqOcQmNX6iQG6BQhef+xG2LLZcBqysngihNKY2WhnbpF7
lB8Af3wjw8zF1WMUqZelRIpI/QHAEnIEyEWc410kmPcZEauPkWhhFk8u0Yr989U5kAaVAF1Y+ZHZ
YIgbCdZSomDSXv/xsN/8dvVlSJLhWVX4weweIqi82aY/VIQD3AHk1ZmyEngsyJ6wS2B2w2MDfChB
LX8vskFS+F/ZEd4RSYFvk76eTBAlxDPuD9H/FiAz2V9LE8YBesADIE7Ygwgn8bex3sA9HndYBGCa
50Xorfn7unhnyfjQXxSciEAcwjgSsPZxLep9aaPzCkysVVd1nr+V+InYmwzr0niAF8VHPHL4a6d9
4+GSWOzCX0kc98cAhUFIskuHtv6u1l7J9z5Jkr6DMsp44BACFpzPfYkPGNWKcfMC9GcyjU4mjdxc
0DyFTdHeizWPahCD/MtExvH3C6jz14Zg5no+veaGHwX2wYBlZV9MJoAvVdXntLBznNEkyESnAvKa
UbYBDrF4c5Jzyv/2w/nBrT5RuBTryv0NujdA+Nt216T5RPvPIfEON+UebmvYcGXHUtSUdfFETlXn
iysSIEqcoBBeBaHtjtMyqV4i/x1nHws7kZPs+osqBvQ7Yfi8It+5uS6SOq4QbgI5NKUYbtvWXILm
nT5vIqMHtIdX6UnC0Ww1IXuz0/zATlnQIcozGAU/STFggjsNx0hm76R06lewPjJZKmg+ubd+/E5x
w2RLI/4/YoaaoxoRzJDbAOwLzaaOk55u/98FRUWOaSts4w/rK7e9FB0276zUbprhZZ0a+Z8WZrN1
csRn5rNqMWWM19JXk03vdKOmMVyc1o9TD4QobP+H9F5DhjuZH0ZGs3GFhzl/0/Du8SHCPpAjgZ5J
XPms6ObDe37H22QbTlGtwQ6aHQujDU0kAs+wwceM0XfDR2n0Q1cHerSIknOp1b17FoLyMcki2lYr
SQq2WNAqaKo/07hcGFcvGoBEh094gFxNSvCy6OOgxUCcodSYC8+d4wSxIqBDSg9kMW0zIdmAevDe
+Ikt2Xl4t+pOED4ZMSiHi6A7gr30Ipkm1FKkNr+jliBIa4wpgg36js7L7uzzhasCoNWT7pgTZIh9
sD3PJSFrnRHqZbrpw1LPnqNOAIaWdXRNplN+F8EbWO0GjCGzMS4MoT0km4QqM0RSG/VOe9Emk4PT
9ZuFNKmxQ5uXU9VtAKTu5dl2YNWD3zirsLH+GxEjSSlMZt9QuGHOD3E2tMcW+3oeO2klrkayeNaW
31ST4okDeECMbj8NiHjt3CiXIRq3lq4BpJxQtsOuZk5EoMdvd6q2BqzAwglKgfvec/w8+cqBkgnI
Ov22PKKOb47yRDa/j02P9I+ULYprh4PAt3ADLnKuQP1o8lFxriu2aeyelWHKUsYKiFUBFjSMyqMg
pWLYxteaRKcPRuyEEv8gsn0GdDRg8LhG6VVuzeRuTDzRPJfmBqsJn9en9+XYRETwupHqcMuh/A5I
FtXLMnEzVKHGQwP1xbx8frMs1EVNjxtjlJAOMTpmJ9ciJ7fCJjyYy+sE7dP5GewyM3fIHl/BGcHp
AcrGQkfmyGRr3NVIzwU+OTt+c2oXnQn3dpzLqprzdTxKGrkph97LEOtXLPu/qTrTAp4dQejOmaxD
UF80ic9+9VEKmCA1Qo5jq/y7+4iJj3p6VmJoBUp6HFHjoBdLlezMhuHcFVYA2llMPuMe3+wRSYk4
MOWe2VKyD32yykEDjuUbV9uTY7S7cd5VXeJO1JK6aGZuP75PomZUN63ZzjnXdB9lYsa+nPnXvLxQ
xWWTVhwa/6K6rw6xXwXWuRigen0Sqe888BBDruiES/HCFW2gd5Qs9rQXuK1ENI6yJio8nwjjA4wr
eBCLHwar/6JPN5WNfUgw4f7M/9b05xc8G8Myy76zYOue66DWBXebRMPhCeb308w0MFy25IzPFLdO
//tuc3d6Twx174Qy4GtNTr2OYE2ewpMuFd0Z+4vz/uLkpnPkY/jIpHs2x7PKorr9YzqGhDOPRQ4v
WgablIPCSrsvMlzgc2ZOYl6Joz6jb7ezT/9jx5fH9guQpG1BF3431+NxYeTf5DpzeCiLjsPBiGzl
2pCVsgC8bXNxopd9zPM58RxXjtD5m0ibthtmPsQlnlg3+PL+qASzxKYLi/OxUggaSJA8hXfMdxsh
XlyaJ0Z5vIem3wR9yM64r6xuiSjknP6cvEeSKu7diuOhZar6EBXdhUsjGO5DD+d0BF0KzrcTMNSU
7Xa+RGM/toVTi3PhE4HIHJyzpMUz2G5zdwh2KXfbwBD0r/eMndZgYkvp3faWVyEQD9z0Czqr8H+H
TN2wf04QnpbRkdqBldpQent9Nw1aoK4ejLkhJr4XO/hulJFdz10825pauANDP7pyC2TZ4J7JdCMI
Pt3yOp/qwfxGULCY52vBfk6RzQ/XStDvmTZhOc49tdBKg420pBxM2ZSII1qtYmVTvGyRbGqpWnSg
J0Q8Yi5uvQAyiHBAYXnL8+WqjBDBip0hpW4B0NH+uM2dthzE7G3qGzuASSGeVeE9eXJe11EfWMSt
zXpEdFa5lFCH5HsgKmLBk1dOsrTJaCwvcUCwWiB0kpW3+g0wZe+E5v6sQ04KLYndXQzUrD/sUVud
ZsNXvepi+lx2gpHw/BnQc0omJTuhxHz6cyFN17Ul1wyJAPZRU7d/Rz+oLJkwhvbEMqPFmAWGO7ti
fyjMvdqyA+7+HlEjxKKTe1InFWM4IE6DkAFVhBOZspGlYhWtFy8fPqkVnVlbbpLqx6xYEJn1wfmB
8LMqeSQpLVX3Dp1i1pefTHQPgqd0fN6pYjwuU/QmVllzAyEGkBhxfrmeKW+Xh2uo/AzQuxKRzQ0G
Q9azH+fB4t4qLY7g12P6sZGrnWzytzLYf8LTXn1OpJyKJunXJQIMszfEzvBN/oB7kbifOj/XEyQm
8rP+9IFwk0YkN4gTESta1Q3GnWTG53OIBV/rtYVN+KxxGGf30hr18Xl7mOGsZkYJtqyFa38HSpVy
jBXaWuOOzBoWQthP5X5Y4WuRQ5Vh+hZ2UHE3CiIDVvtsXE+v8wZfH6TbqOaG18j/ZkPtxVadQVb/
f+VfRU2I6XHY5RfPg7QBELwOrvugV9nGpRAEPp6NK4b0v96mkH3Xj+Sg+z8JZ65d9MgMXarnvAI7
Tak/o7ldzpCQwArqUkJjWLbC3b2B7PVaTvRb//q9Gnisz+5Tur1i6k+fo3NL6NpvZEnDofHlyKVv
VgDfgGpcEj5dWN8vSpg+CK2MqDCHA4ecl+5DvKO7FVD+eMnhGSCio/KJYG1G6SCaBTmkqzlCsQam
XRlkY6wlzu1SYl+Roi3GWfo+OURsZfKqA7mOkS8jKuDHuPIfjgJfgKZXsRN/dPHx//0i/lCD0nMi
ZS9MnKBcITR4HeC5tGqDgNyTmPEMY97hQRDwaJ6Ho7qbugBIIKpXBYNcNPalcGnI6s3N8YE85Cbu
VCzJr/42RKd6tUYVXFGRlbxKx+vJ/lLR/kfaBaNOfHWwoDRHzAyTaS5ESzjxsQZdjcoOER7vhvjX
mYptHGD2Mc3gGhCVdnbdAVa8ICMeRI8xFMJQ9WoJHNN9wdFqxCuqAMTfGiaU6iuH7puLrPcY4t4A
Hci1YemwrvfpYxDLU/9U9fXc0Q/ydtmvgSJ58+uLh6rbUB/ZQ6vrV1CzPcwG5SQxVQIso7i0LC0X
ObqZ3I+TKoZZb3h+ZPxz8rWLuQD+Q7dlxBBiWKoubZfYZzxVSHRjGxp87J+kLfoZlcvVjXjaDQOf
jXudV6S3lrwG26TEuGsToVZOcrF5IxFoUhDykkIgJ7HY9/dPJxe2RwnxMphDZ6bhea30wJLLi50Q
8p+J8iS0cHVdiJ+9c8Jp87hXTxDrTJ30aw4IACENCkJx0/2xlyEHOekBvlcaqlkLFlYA0Id7Q/mU
0v2hQr9p3jADqtiA6FTLPq6PcEcecZoXf24/Ewi9iQJwZukVfUyiJAvS8Yoqj4fRi1YglZgiFxNq
793snW7R4lcfkR4/eCU7Nl+w2Xz7gLjyn8mWNHmZXicZq3fyZ4x+JO6G4TFMrrPih1kcpOf0Q7Yo
zah8MtHEaDR6Eiv3aCIhy+3myA21ziv6rfRRKZ/WgHOyDcvNnvPeLajRVbUDFvfgAcmbGHM5Jts0
aj5Aka2SqAwFViKSSdAn1fRsuVR/fW9rnuLTHzCNhzgDMX1PE/c75EGN2yFLkEdbnFQwJQJHFuTk
/u33TZn9rnr7y2He5uHfdIAtyeoqEjdQUiwPOsviNHI8hqGdVPe/LxXC2g0m7D9uuK0deFB58bO2
u5jqJHZGQ+49psHH4vzMqwuVRcUP0G0PblR+3hwjtcMx9Uk6IaXazfZ1g5rGMSGBp3j9BR90iz2p
FCiZ6RB64PtBfYV9J4woEEK3dQqrfwn8oqik2Uodk9Rhefvh00joCkNdLTO+MsZBokQby0mqNrAQ
BSflwQ55ZuE6skmTLdiowOymm1FoxCm7YS90znk0ID4pvpwluGTDIwW5jL4AWc8vaHfHqMzRSbMz
jUB9VydSpu1AdOD30IjY01NySfiRSWl1b5SYlgxaC4fZv/ipGLHCGQEH2zIwZySWyAUKR0AKZGQB
2bv5SW8ufM3HlU5ZvXhFlN5w9cZSVak69HxrfDAUtAKeLOrw1TF0rSXFNMT3/7POhcfSpl/hlv2B
QdQHfZCavuCN7qEAN7tRlEj2MKxryhIf5Vk7q4S5bv9m23X2Nr1Y6tPcZPCzt+Ykg/ACGP5OEBB7
VASGCtmr35yymWfh7tdoj8MhkMOlWXHJ7hv858IQs2FiXYDRzUzA7qU2IqkbLE8os3bQyEwxLigW
5+klDmf2wREShw1vArJvYBzMQISVU7D5KbnUI978oPL23SZZLlUA5TI6Jx/XIHajGXoVhqos4dw1
KjnAp34KmI4RltgXk1gY1lePUxJtimW9QeiewKQqh3EvTgFzbuMiSXHnE0i1yr0kKRVwp9TdR7FZ
koXVeeUBrLK1+jnAUC9ejKefi7QwBbISgbtduC3oLkX46W8he/1HdNDXHmyaVBScHuixyN7ntTie
aacjGOEqw6ojNG0JOLmJ+966YrYwNxsdQYgpIXFPvrAwFcdHdE6wJUrQYN6I9Fz3UvZxH0zg+CMd
lP9MTXZKYBCOenLg+M92WL1ydmv1d841DSHk2EruyKX1t/dldvfOZRbf6L77IvYhKkP2lmLJ7D1Y
A7mwiuF/UFpoLvRfeHYakWtkBX5gUB1XXoBl8x4ZzPUPquBCb+tjgoG575CwpOKhnseiywOIRgwn
g6zPye7De0rAelltX0B80Ac/V+SRS09bprZmRP2+Hfsdh6xXLsfhv350lkpQkObuScfe37cU7RBj
vt+tMryjtWOdYxT4yesYQKrAV6Q4aHvkJcmtnr1hxbdeOULmTF1nyUydvwCXsGn87s4Ak0/rflyj
GLMxQAnWOoKBOu5Dt7Gm4pN8FYJAAYBsfzhTNIlElsUlj+toFoug5zm/j++mDLAOuVHvnJnxGv58
EbklDGDovat9RcA9njsYwAUkZfHjPrNIVTyaDPIwF9TZYJuBYp+5B5MvmMBa8CegQ08OMCoqqpLC
P6nXFrsvpySKDAVN8CGhEp06q5E9ZRO7qXbHe3IE+OYilsOReRGb9OWiG9O4wBs4pV89+DwiUOEB
2il1kyE1sdZwY0K//d0UQVnljnHFMFuL977l7zg4jypNTa0HNavhoK4gMfjleKGTkgudL09H0gDG
WHSFGHO9PS7R3SL5EnWbR6ZnFKldkeNzI0spi2fQiJf16gKJqb/X5iFsxq6qtLtglZsavyJyjxF5
QtszL5sJ2oIPqhPtjPqu6DEx3uE2CKdLkACj84p0uIWie3l0M5mWiRD27HpxS7E7iiKC2g3ZEyrJ
LbH8h8X36DLCZWZrBtKB3tT3BNEsffdExQDhU+bAG7SF/bcH8NIDdfjbq6BtWs/nk/x7cAc5sjKL
yYJINuC1v8VKimwLVnZF7uvTAV8tpkoMGOPi+PURIOG/vh0qan67ptg2x9e5hFvt4w/sNYmSUAm3
86+Xp3VUep3whx26pkSIg7hWGWG4f8W75mzn/XboV3ws7jJZSm/ghx4S4iB+t51GYz1rmrklOyNa
KEguk8qnGAwlV8Skwo5z/gdRGVu/n7siBvshseCB2igSBQxYoE37POImZmbe3guhgLZkyhYbKgVf
ujnxFnoAvClWcn8zwXkV+hNfmom+fRVoNmB3xBMdxtVXhaFy8xT5SniGNwRjf/SG3d5e8Ue4KPn9
q8Dx82S/LFfVFMiM9PjTUoxFjIUQAiPFFdcE0pjZVBj/xZIulX4r2NFTPljIy9NKeB6du6+xbt6O
U7S+k2Ed+H9k8OmCBjPczL9xXgAEoAekoT9WIIlZ/vQQ3geJSTpav7NcYBjeqG34hS9rgt6RRtnQ
kAsApFSoIBBfuW5msOFRt/6hwSMO40Wga5PGzw2R4WmdROitiQXxIbASIca3v5+aZabV9k6/7vE/
xIv1TlKfB2ZptMNnfa2GqlDDgRSZ/izaTpv9ujWC2owO7gQXp90pNiPmDdmvs4zt92jjOQzxZp2i
Oun36NdVtj1r6ZmnVH7j8Rc7sDveujsB5CgaKRtJrrkVC7sGqPrR4P4uIg0HbU/aXpX7Vl1CrgCl
J/d2oLplh39fBLTfhl1vSRzseYG0SEMoCvNM/fmt0mUng9VXsJhD6ipXyKIUHT3a/50oUo3r2ZiR
KxGy5vNbvmU6qdKcZsxC2/NKuu6IOXfUcXATX/RdpngGycEC+0cZg6XUL5zM/BUJXKMcb6ldBIzU
5kbnY7KgrmsX0dsmDznoJiOf+5KPYArd8+j5cxfwx+rseg1dL3Ug3VeKDvqNr9a2fLtpC5ZjzyjJ
wLJwm9LrCYR322sCCs4fNFK7EtEWvc9iQsP3OW+xXKoiTSMnu8/sl/8zbEyiQ+z9ls28Kmq0iKv5
Cy3SvGtqr8XwpjzO77hZLOWv4rJ/+VE6widJRB7059sioOW5lRSDDoIR0KHnTjb+xf8SXLUfZY4y
rH3K8Lzn8SNetKVZZRcIAk8Y/nUsT8Y5xhu/sSmCIs11UUAFD6FL2/NZXOuRWwtIqtXkq0UhXrpZ
55zMXDMyZ28ymKHsG1NvxbGhc4XWdfHtyXpnR9vXYNuquSRcE5uTf3mIASChl8T1iwisfSIbJota
XttE6rACB2hFwOfcj7BoATyYiACR0YLDsN4PiJwefZ4JOli5UO1wWYbhNQdO3ZdqhJQY9xjs7it8
p7zQpTlPYxUB+xPpggaHu14vKNDr8gkxqoaoAZ+wF4LnnZKw8ujBdh8MfLz9FvXOWX1n07SZjbYL
nyWnp+zMsTfR+UtD1xl5gUXyREN6QsLQ3Ulsnv5OuZu3yHpRFWKCKYddR75k7nlN3I7qbTkODq/j
zQaMsGtm70CNf+s+wc6+9zFPxtnrOx3+DO1z0FuR5XSAp2uADWYwXa5xlJovDJla5N9L0vvMOCnM
Uk9jUEulcvBa0ZwA8mMOU5QIvc0Xn+SLX3b1C8iz6yFltOuGN0hcCDNYkKiQvBf6uHu6MBbUxfVH
SzjlRcj6+rGpeiTuhRBxpAbLAeeDqt+m+eDD/ujVgkoALyT4xTJXXi8Jwy/3kK7CfQhzVz6XpL3c
76bAsOIFmK1Gf85Zu2fKKMlIhUzOgZK9kMClORsxQXO5WBOI6ZM8dRWOIxevoLs0MQAdLQ9Vdk1O
8DwPcsW5hYDBgvRuZLnZnfvnI9IbQsLaM+EYTzkzw65k9exvWgsmixsXA2U70/yOYN3Daf2fDf6Y
b8UStoO0wJBDljeQ4fIznqGS2qorc06UhKvDQZzyn14Cq2XUJmGVgJf8AA6JNL4WRkE92TVoDxUN
B2vbujS7QiNwomeTSrLwjuja7XvlnI9ZL3TCUSXOqMQO6iZAYLIaiHCY78RBHUrqN8MY/1vStzdk
H30GChfJEx8XzNeTLlUyq4CUMoCk8ovcOYpY+YqBkRGL0vM4ezF9xpzAgJBBXes2yN9MtJeQDPiU
Gx9XquYeQSSizBg8sx0qh67Dv48kddcqGyqA3wYAzpe9Rzeol5VGBN07SUK8SGRXxgTPdLLWsqMa
eCIwGIIo3RVKg4vbhnY1BgHiw8OLb7r2kuRdeuQ44NJwxh1ScprlK8bDivd/cO6EDQ2F90XPi44q
rnqk30UP2k3Ak9sBptwG2DI8b/xRkumFzZgdbk6FbAtTGadvoh308GfUmMvU7HaYlL40HzkN2jpj
RitddzRFYr7ynZCwzLKxpkrOs+xBv/tLbNYeRlozeq0ni/BSl8KlpRL9QEk6C0Zf22DRW6o5PYep
H751PN6SQWhI+OAw5dgD36byHJdb+Bt2TA5Us18NobhrfoNh8PpZ9x8SN6dN9QYAnnr4yHWBVQqb
1UMJyJ0/+tXlAoS8jIpsu1Pbc9kXphZ6mtCZ3n9l7rTFsVSavMo4qUoChhSDI1RS+M22Ijjl+SyM
EbSnehGYJll9iVxrrUveyAOsWVZon/yuArSY1AhcuseiquNTU36Q++v2+4yc7jWrTb4dAO3ZMp0t
8XMeXoC7ah/GaMKJJsvJTjoZNo+tgCKXG41DC2vFx+NFczOiDc71KCEa8M6qBW6ZboZ55mdWj3RW
AFbq6B1GBQ18FJRAkh54sOQrPZyr33TOhA9SggEXEoA5Ni4LX6/DyTsgFNBVfC0gkdQEZ2dcz+5T
M9lU4xy59UpujVXLelb9BXMfFeVKYj6V6VoFBVLDGFVNv9zVctQHEyNtgikFdHplZLEuMq3W53l+
u6fcn27AMoRQaTagJIZHdcY+urf+INj41iuGqkRlAiBxmWVqi40eOnYwapeK6xccA9JX+wEuI9v2
D8RvyZmRg3CKeCNLfUtfaEYcTFd6J8WGGJ5B5WfsdjQlWm5rBHV5Sm/jt6UyagOIf09N2GYE1GY0
61LvyY+HY3jqRdeZuV7wsbkfEVVn9wOgREa+xWtbeY393RPjM/sn9oe8Y+Of344nifos46W96XSD
JnT1RTELUzP1AZpBGOuc39QSY4ZdhRkwXWSJDL7sRQznxuZnMDnOjc7zQFYeKXwuU9DTryHrDGOM
kmolVLjx7KhSMsGO7EXudUvSdSyTXMLSKtW0QLGJ/Xzkt+8VhlilCrmxTHiCQ6LY+K80b+E0Su6y
9gpHIsRf2SY88h31O9ZJevvC2cQQcpYdguNPQc/QeEXNnV3Gr+aJ62pgMyrC8IyL0iFgD01CSYds
1MIp78xJyxmh912f111s87PzLoHPu8OuzLFhxRmHXno+m0lrf9p+XbPdh1koEM8OExbMLC2k6swd
O7pi/14pQGJ0ZtOybZUuaUvym0XlHjieDvX2kZSpFj2oasch+vJwbCcdeiRajHurdp6a5hqUOtnB
Ia6b3UfhplHPu4eaJz+oQ74+2gQZ0lsL8CfNbUpMp7HP+ytoQS7J0VmPjbJM22Xru5WOa/w/hbAg
WTfdImOIwlOOpdbYm3LLFvkSm43k+AduSt0VUOBdwJWddqbCivFYi5AlawZQ6rspH7I84zyd1OzE
YQmYJT4Yk4gVLcKtkoZgSMV60lzadKF/yWmFcUCAELggwbkvdUEHHKDnibgdCQ0x4zhOlwCfhzXH
vMOw8VoOsLVfm8xAWVp0FNVYU3KR9HTCOq2905OGs70MnRGFA5hFXzAZEAiz9clAIyUorgUtl33c
VpjS3yJ1F/E7vN9RkJUKNzhr5X5G5psHzmwF88IhCd4B9ga44gKRMRTPdueA2zFWlkTxq0uKodzc
jKw22Oj4gK0olaCqAa8eUfnVeCu29q+M3Ph0H8Nj4u57XoCi5OJ7kOYi0IyoigLDl6WZA98HiFVw
UBnIwfE5qZZF39inix2ATUxlRK8hkLHOUexL0hcI76xBvgpN54zVnqUqtjPdeldaSVHVYVmVkKI0
9uiEwZ2VcMGCi9DF8FdirmKCoSprvSq55g9RvoNatZJBkZCcFeNZArJjlW6SMGthzHIeyKnGPvDc
5t4+6EA1pAocoYGNG+5NJO0u4k0nii3Y8A5JDjKW4ly7fIoX2cnDbQLaBBSsZW5A0xrnO4HhazkK
irbEs/YXnBcWmd9bRkI7A7xWWueHiq8oALGIKlgUD9LaoEBhYmPr6ZLZ0bXFiVpV9lIob7cijeQp
OQvfJ4WqBT9uH5IMty7npWfrSqQT25Lsd/QL6hBZ6u3EgS9D5q+G/pJs8dKy54W8OoNamVmbF+1u
eDW97Y9PhA59b6Fhb0NagKS/Z1mzfUGDko7b+/UQ7/qfRbT5OB+Q7yq5jFUj3UfP5iACAWlO6SjT
pZfg3w/PFhKA5OcUG+G5Ro9WNxQ4K5GrLdC4PDgRSN2kWtGMJxDRSFT+y7tdq5g1zhWlER4S+pHn
/85vG/Di9JxkD0Ms5TCUNgrHw0nGz4reggWlOPQ2RVB2vBoVG/q0KOPjv/uiE4LV5sPLbP/po9+k
pi2asOj3KWjWSzZLvdeZwCr96xJJc86f/EWDPKhJ5KO7K9ewqp0h6RwjuPWBLs0cAsQkxgbRxp0u
62eXLczs/xUol30G/gdPOTFAijv0UQiHiP11VNFpHc8KWuU89UDIzGoiV+PzLtsGYzgHrIWznV9K
11VbwYmIm9GmCvgHRK0TPP19PuG8rQcQ56DUMcvwrrYCkC6cm6NrpsUdvsZZ4bQxu+7ERWWldl+6
Zz1YoqfcOd1E3Bc/RX5Dn2kOAOW5dIX2qIjXvP8MldCpWmXhaylNwxRlIv/K0MC8UNRLE2az+Ap+
t7uPjJVcbxfC3aJAk9tskdogCHUGCoBypMzJEzTHaVYHJvmCfdJcAPOPHk+La/d0VST6vW1XHO81
9YCgijFprtNU7tcC6HaVJOZhEI+NL6NqEbEWSZ5ekPZqlZe/rw1SNkXyeFBBK6C5X9WlF+bSIjk2
f+ITbPCmy+TUX2mS5VCKEbtjTJsJtb3V2dJu38Ug4hFKeFz8Yn8zy8yrlC7OGoNQdR/4qqKKrhTe
VCdII04lgG00c93IpHN687VcTjrOxnuOrIKOzYy5miHdE1mG76inUSt9AXWsttRI7leVtr/P5XhU
vlJdeQw9UJZMYMUng1OzINMLvxZFpWq2/JnAJfYEqo+aKgl3svpAo0Db7oPu4IRGXbow/OFsT/m6
4oBjoEfYIUs3WFBdyY+HayBUGfkz3cw5chD6ZTJzm5Vrb5jPns9XlR2unbdsk7/awmJm/XJE06YA
2h4Wa5ePz7MNZi0DwcvyFCHhPQuJdSCrAmDLOdyz9VpQCN8q6ZCEdrgpGGEUAH8XcJcY5aLdzlXj
PAnD4EoxhDjdws5RRenjGV9nwDijYii1QlnKN4OVhMBYgeFDnmmAxz/8SMPnQhYdVQxquae+oRCA
5yYK2ktzRXDGlSjNHSe2WygWcAa+VqCOuvefmQBm3T6I/9MwvZPxuAH0XtQ71+OffE8lJAp3sWI2
z5+HbvJTLXOeX/R2MqJkOfuEiZsD6NuQGjaP7MpQ1+sRo9iN2R/0TetxvCx5erbZyZFfQmv4PgfD
ZJf+FS7jMQK7W1AOilDGQ5MRBFAfKi2gFCBjO2H2PVjhl796ljxdzxJwsucZvEyRlCuQ0lqACxFu
VUxUeQNVD/d2t1K6S7RF1d0zMKUko2kfiPHoEAw/w/YS+0Hv2WclPtgf7vKQZLxsZLt4LJx3O9Lc
0pcSZWXFXrq6Z8QdNBB+HkDxUkxlEzMJPIcJ/cYU8tHhF5nEnfg1eacwC41eQvBZu2iEGhQiEe4b
pYEV2FKeY7DCzF2E7b4hQHvc9UH2XtVk6ShjZ8rYT8aRorPvfZ+nHQAR51GJCtNn7LL7wPlqYNTv
w4NCMtpShm+M1Eu5VhdU6tUvKtOpm+uWzOQy4DGsJ/qUQoEMWjVhmi+OwuoSa8ThiwAsRplbG8h3
3ORbrYEstxGQC4JlJnL9QfSmawkB2aO/ymaTCPo9R9UzfNDE8MSY8Ntnoiij+jd3bzTyOEtXRdnP
WNDrQ5W87DWVctIblfLkoM+rQ9MR6Ae8KMgtiLel0+71O/8iJMTJ8ofCuZrznhzbIFqeBFyJZjup
zv0hpGNBYUBbBzabEBrm/mocvB49nClvk7lyWcYhTYVcvj1Q30VUSHNFmJju7fSkr5Li8MvIZMwp
ElIMLQlcRrnlo9dAEuwSGxUa/bC9xpUesGcpn3czApO/O8nAkfEpiEQ3s1aV3Ep+k6f5t7MUzRue
VRK/VCS//FgrPXS5RPfA21+o0cHkukO1dxWwWdK87M6dEA0u1qRcLbKu6vWfI+KqxlhQFNDY6RF3
NEUoPa8tyJ66CD5FHwzsISfuf20aTPCAN+KLuMvKQe5CR/3l/whOnfNYEywNBBExjUXZEBs8XgYB
zbAjQfEI04BHrUYFfLF8E/dYbgZ1BeC0cswtwz6xlVS7MMMHZs01JO1O3bkin1m5WZCgnX/SWKWW
oc4rOgtlYEW4BOhWE75/6Kw9+uZU9uYMQN9RuUoEEC5FFLGwX6V/R9V6BRNjaWFIIXviZoxvy4IM
+dVn50zGBO28ne7GA+Rva76SOne/7kFuOfBl4r1gSmdrJaFdNK2yQ16elXaZVY3x2cO4AqepyRUr
N3O+hSYtSRqTubXxNs/BT7L3iPwT09W51Xu0AgPX2dR4z2BzpPNItM403+9cuMSKrcKjwRfm0I3z
u2mafZNxAAqh+X1G+Lzq++TxKu5keMKh6Dn8wJaiam7NQmfUe/bfuUvsI1Ibu0uZnYPtVqW5Gjaz
bAuyvRCNAp7ayACBtVDvCo3qjNerAaZCBIGUNs2zM8nNqJqvsR3hIRfDjXmGN+to3DLJAv0du6/q
hG+rT8GZS0fcBVdnwbAv58XyWkdoo+55+NCV6h7R57JrfDy4nsmYwjYId+js7aN+aAYijs3bi0Ji
Jw7ntKvJBLPerpcZkUKoAHrducOPQ7p/u+KjG9aExY+Xz5e0PIbw9zBvm8hezGyB7cm3QFH8XyKZ
oBeA+rArGRzBtqOV0cAYOdM8M7k7v19H2wpuFklBahKKIqsJ4tjsulsvK1OUPu2VIJEZyw/mXK2u
lW/9pKbPcedZnesGM1gHoAjIa1givdv0pI2f7Q6ClykrFdeIRUpgXSYyULWddpb1WhP6dZDBsJPP
fPJz1OZj2b3pDlJWlxiDwUsUSbDHTRGUW43hskK0cLgbcrPzSodp/QxmfIkSVpbgDdWsiUAbgUav
gvFykpgxWk//sEVQ+A1E6JxVHKC5WgdAULtlfX4/5Po+B9OL8iKsJ6dBIe5U5P565hCy3d2ZgB00
SiQdnzYfdlv+OEZYPMNnYhcSS12J3u5X8jRFQVeLn107M2Azx4h/rhkrNoZ1MZmlQ3Aek/LvdN59
Eif1madCf0WkFOlkDW2XmOZI8ikvuci6H5usbNKtSUBdrjb4g10YSMwyoXpdKox/hRZ6EO7egurk
R4HlREFarf8lbhrf7JFOfEvoFS8TmAw0heM+PYjNG1B83hKyroii8iE3nLDguSGftpZVLgAYtGr1
vWaSOHDFKOuLyOTLndmFnUmSRv3EUGuYIoL4ygiztcMT3I6FjluaH6Of0KSE7hT/qZWAlg1rM01l
sC3/2zXjtLcAG6CWm/AKNJgGzMdXycz0DCVdSpfepfeKa6U8IWHPzHKtwJZenp1wnfukg7U4thVt
AIusVgSg5zaV9/y9Mhv2EpzR+ZBAYrpuHsXJ4o/IXiQiGUviexsBKmgKxBc4vDmYo9es0VLIvwhb
hArFM3fRAytFkm0jMv4Hryj+SqgK78NhFIiK42tWMWAM1ajQCx8Z0MM51Ja07sOlOE7g0mPjTNwR
Gc8QXsb/cxehBE6veUB5TX35Q9MXDPAh5pgVYaLgP/8QstjTz2MqBFR05eGksUZ8fY7JyVJQT0II
wHvTiW9hty0oBgpY+r9zq8xuKyezGXDQHu+qwd+7gAWkLDjmb5xc89+kw4jwGo5uQe9dwCnpmWva
n/PPe4MUqReC7e8hGe8llMdAZCHUB/ZPBVikk09DvgYQXvxdv4Nt4hBSe2z35e+z9MNug3r1eHmX
W9WqxUP86YPVw5UdMke7ZaKhMkHMinF9r4dDoO1OXozy1R9WsxjolQNoHrx+hDmsVUWGGyRFpu6N
OnckJvJ7m8Lq46u3jrspWbhPDhE3AO3f+Z7fVS8ak8bfLNdJBXoaxEjcEUjZ6odEbg9Sz4AX1nuT
I219emkTxHetvtQ2TZldZ5sLJmZU+iciED6xIhDWfHiIcQr9wRtyPvgOgRZqH7uyXgILR63BBPbC
UdpeBKJAIirN6Fe4kC1vaP5Fxy8d1nHBxFtpsbCSo+gZgq8E6oDOdf4W2fv50/wseBsmdwfOa3oe
cYZLosljwtQVknDy9Ahc9Ju2/Jt06y24/t8zwQWLG+2Z5LtcNQ6PfHgmhQDc4tfmDmDRJoYCF9gH
dauHqNHAb02hN3yu8uVlrLXqdRHNN5PXiCDKnTwCy66qSs8Ygnbp2kWfdT2Noi+Im5/nGrKJCC06
UC1uiXQVxtpJH99xfgp7mmBDMk8I047UqcuSa0bhEYIdtOjCLCbPaogPPwW92zYtuekoNkqgEOfb
YxI6LkGPrv8WLrcOi3qYrtf7i78jVhpnv5jUnLEBb1cFxK7xjuMp/53sG/kL4+wcF1zNVqpTjvO5
MMe4OdNFC6ohyhBhv7Zgr+xJoXkv7YKheP/bSSoYNv9jisfxQQmLg4rs+E9A/Ejbaiyx8mD8HHJI
ej9wonfP/+KGpUpOsICtxV5iiCsa91KWaWpZAP7y2s3KnBTtQRFXeSRbQkqa6GEHIn6CrmCTBgBT
9PcBwm3zEOvLidX3E0dN3mcWX5jEa9BGdWDtfFqQMSA30/aPxJ3HkcvZpUtspLkAEXG6OVGZJRN1
26LYKKS0m948z0FLWIvTQvvwDiKk6nubhDLZMs6UcWCRvfF4V2bE4wHN4+WirMNITSefnnT7eGYx
eQWc24imkkaaM0hb0fVY5k4LHrXlWLCMr/xAm5UC6rABTEh6iwehu5eGCRCLj0imEur00TebH3L5
YfafkBpDDPzOUSyDNKxrYF0iigFsY2HUBkYcPpKN6/f8UfFAzD8bfn8wigqe8QaULOgtOQxW1YAK
4Il5f7Vk37wW/Gh2stZ0vFy1iT5MlKWgABYu5voi8aBoxkIxJznyqK8/xa5s2sG/Vdbf4YWe4Q7k
YWAkuqwg0PdZZ4lHenRE3JnLl6vZqDu6qzS/fxeluy6EcdsCCCxXYdpHCLQZxn8hRSObbdPDibQT
Kccbx8OkiZJBf0bRDrQdt5rS5fgT64aX4Js72gexGodRlLfg8q+m9rxkUhoCB9WyKEPCGnYZeF3z
Qbqxa6ZmSQKq5DTW8EoDhHb5g3yykyafBrK+H6rXFoqJHLwfgiOPbp35c/670khKSfizep4ySTEG
G47VK5PxLS8I8M4g6ZPyf/VVkNkusNzYSnxmHNMp7f1h1fMTBf5O3Bn/UdVGuJxBqR34L8JgQ4ZS
cCyM11p1hSY2yQjAnUf6qO7LRILmtsR2BJ14FTQU8NrleeI8wlmYp4+s40wkPFkaNeyYIfaL6Bbn
ANCst9rhgfUyDdw5UW75uBH9VKQPZ4w6juA1bDZeNCbrVlTdAxHXlXlVQSpEt0s+JXr6fWuFlXAr
n8uFkS9BQTzd6OW+Ghae/f74/RFJiJw4QWcPqD0ctnfazpWOQlUrqDfdlbkr9YEX0w2Urb3VGzj1
DcXXteo3IwouWhgEB21jrSYVI7ODxy9hovwvvEKhuHTHPZn80k/4LxWyzJTK1pPBFl/m76Q4O1Oq
ANjR3MFSxhJ5DMI3Csd/CTyyRYrY+FeDW+2N/FyOw+Fv1EfjSypEbp6y9pb3la8qTDZ0RAw/N2P3
Ryfz6enV4KnplZ0Ei4Wfn5fAREUQacPm9u5qSn8Q44lKA1cNRyPZ/D3Go71JRpyDXzfHupnr2V2V
arTebjvyKC8BF1GqgqW7wdCmducW/MqTW5K93YDpeBf3yVo1PxxsljmYTU5wzsuNoPswezQ6aw3U
ZzxVRztYJZ406xz1PMr1N2Sk6r0zb259yYHlsPnekFj4wELg3uAGAvISYQmxk4SL6ToAvJyJ31rw
UosXwAb6ThPegDxira8xTLtlTl4wXFq2hNeWtrQ0DnZf+S9Ls2E9NSuxnLSdVSNDnnZNdBE1v03z
ZMvmvxIe+IJFSDk05KMHL6MCsBtRxMiYXBZQDY6CSNJ76mmqPgAPkYICZOxqTVaSJDG4nmJGFd3/
uL7PT1Jxsws0WwUgzXlm5Wfn8JF8Igb0938rm4L9QZ4nGPDATEb32vXTyAP5xMElheY+AckuSCdM
th8KVd7wyTyl7Sbw16cI8G/4HFU9pnjUrOFjrETTs+5orPNobEFmepJ0vQm6B8RKSRmXzRLRCGFW
7uUidfXMB/fcOpbUkWSHmmbNZzGs58zAQ4X1lZR/guZPF02B36HqwUXJqNCBJJt8a6jc5YuVe9EJ
lTBk8xI3Wp2f4vOZwML30x4XyRxKTQK1KOmSO07w0mtXH/1FvoTxYQw3PCli992x96c7/rQ75l+M
rsCZbKp2Smf6mcJt2I8zzRiKxgWQFQHVde6Az3nCVkkjYUxoR0W4xLCsIGXckftAT8q0mDS1MzKH
XGcazK6M1oYAhupdSpuKopT1AXCqoNkULgHt8yYpKPmAYyDIv/ZuNh65NNtDK2vXf31ei7ZYEFgq
CHs3eIxT/ALejSZPhXTgKIkfqg76fwxTfn3c5iAOSPWMSVDO10D32+mlGYlWa8GZ5vN67HWE02+2
fsawdaCF9mJGrsL0UQg7fZZLf2Oa7HenTCH35pg//+PhE8klHRK7/9MaYjyo3W8gPWQK1SWjWDtV
VABNEzNQefoo3OBKh7AMtaD/KlbGyYLjt/DMqcSOxVRSl0RP2u8z81WAGDL5QeQjaaTJNhagPATi
ATN4jFo/TKvP0R00QwTDRri1ZhOVxUeP/bclU+Yj1hXe4huNo5wM1REVdgWyBCxMgb+5I4EYj9c7
FQmBklzIuykHdY9QMHM6JuRMQP8TRIPVJjEMzKj1KkDfmF3VcUi+MrhBwB87ubAevmki58+o+nkJ
vW51xs4pYbRthtS8BslbZLOIcqSwhr1/tUJjW4ebMR2rRERYnzR8++9+N30SwyF8116h8FMd7rK2
O84dBzUxdrjria+LZRKU5vln5UjX1gHq/HkRIQZ/p+wQqadWQZeQNRLe5vJ9JHnkI1BQogDxgk6k
EGo8hEKHQ6Vx9u7Js5LSLdhjoPZMShWc9fmIEncR/XKXtne1P98g1n6ZQB2ZwEHyEicptA6dVwO8
Trt8yc+RHI3t18sZVxIjTDXpOZRM74FY6UXRC3te30FkLG3Rt1F1VkaexZyRNK5wYMdRTBSRgrX0
y5mXw02msXQOpG0bzslYsA9PR6aO29BgVW1qbcK0+LVQjPKJz2hxsi5QwvnmPypG9Is0maujQ8MX
akANcvjJdRBqYklLcUMriFzVzrPYZHSC+6gKj6CneBU6brZNLmM4fdJ52PPrd89lOXeJCfbRCG8i
cCIBop3xB5xUJiQ64WsQDQSBT4lg7VwNG6JPsWsQ61UOlgKhE2jKdwEUS/cYqw7W5dreKc2Q9ovx
xp/MNMbVd/D/KDSTaz+TiKGl9Zog44uxetqG8srXTJEM9jwq/pyq2DBQJzgpVvmqEGL9sbBrHVyR
WhHSiC/HUdwrKKjfaGba6qIz9FYWmk0W1AyWmG3K79e9KpkybCTVs+MXNQxPpkxUXceg/VaHFH1J
PIKyBZI5LJUbPGLmf5yhhz58ZdGjZjQeXIB5Og2yEZL9i3MieoZP5GX+O2xW2F2nU3+p7XFTYsIO
TqZq6hfLIQqiviSvH2J/TQsUXCl2k3bZkDGiH80Qju+bMC54nU3tJcPAmFhJu60Uk9X0uSnIBprI
KOgfQ5JSX5qNi2Jk+0aOVgsXQB0hUEH6m3mdGnhJrzZyLpPT7o/XeKb9rwdCPEVKkrwyQrYI81Cv
0zjVsks8SD2ud87BPYS3OiZijLuhLMbUccOZnicooEefww1GCauLcP6T+KGpgYiOieGZzCLB8aqb
0TkwfVbC8wXeepkK7JXiyLeYsOWN8AWeanI+ifGza/RYZ6c9RJiLv2XwbRLYMkkOV4mazuTJRmsq
EweQVCs6DXl1AtEaQ3bZqnmsHk+EmLp7SPRPLDuWcq3uqoD3uNdJR7LzTcp+2cE1em1bD+zBiGkB
OguD+G4yKu60V1n+NEdRf1/6J+SP5Hb3a0t/tyKK6f+JixI26KuomY+rtMRBT6jmlSo0BKPgJnrw
VxzTtQ/g/RQOtP8f5DkaWi1EwW678r+TmecBpK0A9aP/DN8q5kD9i/LHHvZbWu+X3mw5GA62OEzK
7+fizkZjTO5D0pAlG5sBS8z4E9Nh6Tp8xNqg4PtMbpGm80ImXbeCXa8uBn44tpYGa6LaChwA0GVI
EKjEeYn6SHTghW7QNx7x4WKARScyOFIaKXPcTHVUR0p13I/h6HGK3S26GJyPRL5wDy2H9DupiqTI
M1AnfnZPZ1ldQqyOHS+63LMFHeyo9sl3Z8rHvFdPV/nGFShUyQDnIJwAjw+AIvemUslfj8gp4Z24
kXcsob7H86fuoiuO6WL5Bz+pjR+gHgE4NsAxBjQ9JEDoZb+BYezIR/k15xj3oeKx9p2zhIkvp9JK
OnBfcV5R7I8off0rDmjP0VNCTnDxOy4WjYxGiBUWCk8gipXdO+K9c50LP/QLG9YMtK0PkxwJsKiM
q1T1xYiDBXuvsHS+qK+RLMIct0pS2ES8A0JzeLrIvNMuCBKblqunsTao/PoK9+y47hRP77wFLpNt
AcIE4BehHozUWlOe5c4pW3mdYMHBmGldl5Lww1Wb7FwJjuWsZNw7Vd82hGPKmEpaCe5Xf5ieQ62p
SN8mM9r9sEGZgPBA113l6wQncfceEZhwUIedImRWHdYP3E2P4Rfe3dqdHmXJ/OaUSO6HjQwcnEe4
SKKgDsSmI3JG9EAZ71IaOQgAf4NF9OCF1SuvOLsxk2uNKVvoqqdxgpLg9Hm+FwQWJZq7etwL/smx
eQRgIYjH+4EEJbdAmhC6tE034Lgbe1Qx+knTASord9YNSUmK46uO+uKjVDfwT/LYY2Pg0F+cDOLl
XD1aCD6c0jpPGCRP1saD1KodVuP/w9/Vjcs/WwNp9gUiP2BEyoq7o+5TMmuP8i8T80f0saiee7eS
Ko9JoMARzGbwV7J1QNBHj8yX8ahzZKrkZF9C7SC0KzHuzjVAD19oQ5uhKgR9UEqM71apoPioh6KG
ZzV9K62Dz8BQM4OekStJM8tHqrCLcoSfPqz9lHM7u5dy9+9WL/muXVUYw+3K/HKptMsn/zHArriH
6o/2sEqneunbtREfsuI3mpmyzwdLWc6q3MJZRAf3ayGARLapkjqSD8Hud4MAzd1HlIl24uIdHq5V
iCgUCWWdStVY+CnvLkxz+q0WQmq1ioh4Yz8lWut+aEU06EM5eeAsuIETn8sU7FHQp9BeE/JAo9VH
iTPrGcZiM5UpIdCqQqJclHaYG85dnGBtAlWsWnhWTIzwIhVs5HwqakLcgB53hCPsrbx1XvHVUOJk
S7wWyu4Gtfionn6/rfklcsfPAf8y74xyFCrC0sUrLFC/qef0rPSnN9bNSYEN3k+/bR7lDswCi1g+
BAU9UU/xwky1vdInrP/pPVk8/OVP6drBvaqO/7HNH8DMMJRyGF3LVQWTmFecF+sZd8FLt4RJFx1L
dUk+Fuoin/NCevuL5sAik0pC7kbGZmkl6M1HKwCGgGgPswJ1LHYVVDWM+vEkKnD+S33T+VXcm6eG
RqqJCjWzrHOragD6+6FGuumT0bepJn7UYCU0z80HUcMRAaYPsTd72x8b4+rfIXhlkavQOSzsOv8p
bb4ZnNjBar8OuT9m2nf7cs/lmKGyLeJzyfDPb0bgjweHoR+n28PLzO2RjuGqS67qKdocYM2zMxAk
pU6ZjkMPW+RO7jEQuPth9kIdjTuAgDYkEl/cpjww61wtxkzC7o2EJfOW/xMPHLwJBXDPVmyTHB7T
F1K6ZGg9oMb1PbkM7dGq+V2aeS9G7Kk9yeWDNsoWYuVadREdyFh4DBvTW9VKt1Ymxeb17fXHcB61
ycrJEpzpHj5mJbd4mXj4qfoeSok6VWH3D8Fncky+SV7X5Qt2G/ZIUPyiGs/jBeUmI6guXFzfOLgy
ZLpBkdsBi8v20GNUzSYV5Q1mmLiZ6POmkHWMBzy2o0QPM+Siqzup3CiQ4YWPMaP1qZuCTKyDkJgH
UIKHQbciNDnbF2kv8uFVkTcUWjhbE6aYguM0vNF6CycEZSKICpBZ88ufN9EXE+Bxt8QklUpYeLAd
7V7lRR32Bs6ERJq+QWUFNVn1v+rHaL0OcmJHcM8rjhyKWMFhkpXyZ0e/VCdpZ5img06LIDNe2zqk
ue9/N5f4R7FFd/736qOj2qCioUUMhen6wdH7aEg60q2C5yoiAHKZoldgBFMIxkolmFy0PPOyL04A
+txGQm+tBUm7ZPmTnXfhuWWikJ8rpEcbJji8dPLhyv0ZCHnfY4Oty5tNnxrnOz7sioxrmQMFO2uT
n2uSU/CmXfwHbCg4PLlucYqe2IC639yWi5NhKvBpiJYTJqjm5KH59HHz+kQSJHVgTqWuWSx6FQE3
+izlaF92pgssFh5Ui2UaEXRmWm9wf2YNp4zuyrQ927GbFBOFaMLEnG7SyrXswfETlfaE86EC+fqR
HLzM3NWZ9TipEm2xgk/kb8w4IhOFUt3RblkxXzPUmKweKsG5loQ/aHlbJH6pnFBMPXgVZxhcrXZV
AsR44PswUZB7DTAmwNJDq36GRzR0i8qSVHVzPkD8QCi5VqvBUtWmG5MS0ArAD1jVZX646LwnCgnz
JF1rR0KXP204uV7nNBlYTDutmi2RQ8dFMDCQl5qSk3PAzXYseS2ZiSeJIXJD8KzRG7QULvbz1QVl
qUBosWNwBiDcui1xqty0XELpPCCsNcxtVGlib0NpDe8TSKjBs4+/I/pKXI3ffEDIzZaQyX9CSq5m
RXthtG89jlg5/QU6miUxs5clV+zAFD3TomDrFQb7jpmMyhm1OHeAhsWe5D3x0zOJk9h6YEp/9Hag
lTflNmvcRSlt27IJLSWEHQEciIjAkSK0fkCzUQx1skUfVAyGbFMBEjeeM/fATjwKBwlwpLKJgzBT
B7bQHUQPAZPCba6hzVqTfvfdDkAXXd/mTDu+HhPe90/k0TbqXX5H7WjFXHnnIBHuCYY6nRAwCLl4
yhmtO1i7uKHdI1eGbFC0vNZPxLO5L64BwCkD5EkXJcjWOkS74UsV4GqaQmu7X+G8OGdGI2Q9D8N0
gMjjK/3BRFkcd6DKt1wHv5Ei+NGVoFvia0pnLo/1X+IYr3Z81dPha4f5pauwSrIErOO1UDnqYuFO
qL7RWlsEr8hwBCBxOa3WDqmuW1KW8J+TKQvK5bGKgz38XLgcJ5HNGZElkBSgNiVSEeg5MKhlxFXS
mIIyYrQ6EgXFxapV2OQElZ2CUgc6gbmREW2VDeZtE9y7IIChdY6Km4gHqtTc3sUup5FyhebYvvzw
ORPXBtyhUUKI+cxE/FSPotZqD2BFMsfkX/tcQGc83etUmjELvnt1qMKoPDzi/mQPCL+80OPFjHOW
+0lAlRnWtGbqW7u7KunXNSIJgztcxNHXfhy5tn5N8/Qjvzb/u8a+GlGOE+YKbME+kKgvrjH9IcVk
wi03NOdArJ7V6AnjjPKKKYaobwGbd6Psa5DJqmfE4HnLV5IYZ8h8xRV9S/wXSlEfbQB6gOsc44Bm
nNifke1UOVafuQp2mwXntInvgsQhJiLFUZeIvtracZbKlE5JM/pX0zjSvmMLIiQsnhhD9W6GVJGT
rAUOYzbUrlpb4npbzYWLpDicQKHtIvKn8Qmic62Z9FN/BWv4o/iG76OXzmFkpZy89Sa6yTCe0m7l
k5zhDggtWEkSX8PlR3CvcrB3HhCUx/vOdPVXHY2necYpYzNnnc2v3gpii8ignE5ceZIhmR+U0o6R
Dd1oFpLCYIrqK3gyni0itT1myRzbGci3dOltod/p+yFDB4PBsCPJiwi9vtCzeEdwGD/bwr3VbIyE
dRtXPSBAdt5XqSnCkA6WHc46P3ijbI1afOOOUkvyDjCYUJrYpLrhmsnSM8xalrZzyFKUyqpSE71S
V2E0yhGb92ljoxjoTeIEVuv5+eU1FRdu/5q8XV1CeDHZnQYevriWjXjDNjxFRxg/Vz4id+KKRIlP
HY29OwGVdRKkE/r/vh6qbPkWGFucavkmd/zfwnwmeHcet89DxA4+3wMKg47tC0WF3mlnJStcOd97
cVdJGdEnjbCwkKu8JgRZyhnpqQH65eZyUMbvJKA5CLY6yvZtT1OHFYXxUqdwFCkKAnbfCv4Zj4p9
VAfLD/crBGrtDO0QLC97ZZpj9kpzqzU13jJZNVkyR2BV00QZiEi0Cg+b3KbBPiBExlAMIUmNse0c
JoHFpxRHMiaxCHbc/6pgCwqIZuVq+0cpFWnqCArtsqO9fpqQ3YFX+pkEX9Vf9KMXEWCdCsJ8jjFz
VdcXQv7gaaWQON2RLNRFyeDnlVjrSCO2PGXP88mjz7FTFrpI5eIEB33Ey8I89z2yzdlj+7sgEy88
3dMVTw2vrV1/fnjEPToe92lyzQAjHwdfzn6foZcotQpK7jxNHh/LaJDbKG5jVkoJxVJLbOgl4Ckj
znu6cMh6QJ95BQkVckOS8Iz740NFyLFzwgSlPfezR/QDCRfhURCs+XXGfufD/7q+T+ws0YMJOzrp
FSh3XuLQzw9/ctv7oYOsoOepJtt4lwhJs15wJzgjp32joP0c72NwiRyryzKO9AxEw3R/roJy8dJB
Ppv/H24+aGrDlAyQ6Fd1J9c3jq9XfKa1sO56WNnfn/MflKfJ0ofcPXlpcmqncB/i6tN7FRr7xxPn
6o5/bVWJpXhZusl7ZwRi4t6e+MAO6Zng5wZI85gQTg8ABZlANf4xbzNuFcQ5ME03jTAZomG+nAB7
ExjAXRfSnV1wIz58ENiQVWTEMVMDDjNFjUuyE9E/boDwsuxmpKUky7cjDDr3Q+hHh1uTDIEROfXX
QBUea+EILLoXUzbAjO2GlwhtpQXMcJBn4Qx6g26sMJMOUsfUfN742Bm5u4YVv8qc7MbgDfox/KgZ
tMs1Bhua8mdH+X2Fvv9W7VcQS7LHylegwbBkYfBRXDjjfuU8Eg+4itdYsBXs0tDVzZg+jMDwLGV/
1SC1pJL3LsdXbszfAvnFff9DBE0r+u8fluDCUOpDUX8FHEoJadDkxQwnyEwCEKq/InO8hvu9AR5j
LRyIGutD9QNemOmhkMi3cjw+b1+k+uGWDj0PdHC89vmcDuSt2fxBHyCMjyvlpMgnrJ7QsThwKYuU
/VirxwXjVrthu66kuSi/CT3k4NfhXSuQ9Enob6VzxE1ek7JqBgkxAUh6xMcBgVBuEkTdhY6fceNK
zg7T6mD6YqptXiqMyxo+/PEa5gWNX/Z3l7kFarsr59rcHmBvZXRSnKY7rFRt6bVJYsWY0lOr1Z4l
r4VNx6MGaCd063WfYBNY8pO2jQhq8U5LueND24lhCU8VNl0002MwoLsiIMjTHpbDJHQl/j9yHK9y
KNMbi/IqYCd9MbdFgafbAgLoHFHqZrWqT6Kx9CInGeKF37rcoOK5u+ZYQ5lSVh5G0qE6IZeW0W0U
jnlcFv4ixoK6gKpBYIFl46aBkV8zytCLcW9fUw3WLZeoUoYqKfG+Txx2FeUyYfvdWBHN9l8zibH4
UAd8xLq5Gun7mLb1w0tVQZuEpw96MPMe7hO83R78sBy71mqGH6RXYdRDZXeKMGmBS4LwyKuWwNA8
mFnarCwgrciQNJljLQXg37hKhbCNMoTB6Xc2WLhU0z+nzijFlUtCEFlT2uUfY1NPYNVaLaHliB5Q
F9OdZblHB7mP11E7f4e/I8PLJEc4nWiTigo2B6pipB7cvhx081CXxC5kIozCjD5fn9kcqSeT7RJ/
hdHps8AELe1bKh6iCGXph6VajZa3al+Ltd1qJ8dWVRS5bWfgoPimv9p801tqYXqjOWVnhJ/fTzR9
i1SFdMYTlF9vevvjKRdxSo5Hz/4FK8li/7dg/3zc4OH20eekzEHuzD9mUGSp90WDVUWZbWsEej7n
yHs82AT3Uh8BHfwKSV0exsf81vvxo4ogthmM6RQOiQI4SNx1LN1jMSCTtpOUn0aQ0vCNZmznB8he
2Zia8azNOUkJJLL7+j+eTxe+SJG5iQMSNWnCM/pbAWtIhkrMyDq6Gmr5JLCAhe9srRAaUQuCi+ny
/CavD7aO4Pb9K67hPqd94sJ0Njjq7VrBGRWTZ/d4f9C5iUH0l+C+Q0JtE6nUFwz4U8WXr2wcTkZW
JNLZr2WvnFfg80dKS5H2Hl+8dxpRyKTrKPc88N688fFTabWSLB3lQySDXJJvVeM6fAWgrej7g0Fa
znOtdQLhZg+o77ZJJ4zcOwqFLDeBBZp+JKAnjC65RHvkXs9kS3RYgj8JI5Ah4NdTKCxUhwD8Eboc
y/nmIqdE7OQuAIE0DqbSqgZB/WEFqg8UDF6ID2yPGZIlSjNZ3aG3TmdUQT7zkAHH0v8B614J2P/x
OBVJ0ZsV6DpWvGyhn7mL6RhIBVjn5ckL87FrI2gLCRWT8+Y7kWSG9FPJNdkmf4Q75U3JcaLz87au
32YUnm1/M4Sb8nLAiHPvLWRQ66mAzGoEwk+cDRThcYRUlBqDWmpf8IdjEVFn1kVl6mfBhr27sFrk
bf3umPQrQA6MV/0wG4AkHGZAGxKctVK8TH6yCeu051vqmAQ1+G4YrdlbAuoxfXHbepQmR1UZZ10n
+V7NZ7gZMZJPvi8BSYuwF868TzflTUVfZsuO4cwe3ZrnpfQ3aA0FqiPGId55feKFzgENF3fxtGq2
3fF//9kXPkw8FTPCa0cTVxLsvMdg6JHoELe7bJI6+bHLK/aK/3Yg/AfcoMG55h4aySRWxbNbZaeO
kXvoZfQf3fl7PWSEKv71HlHr0nhL+9dNpFCsIvuBMhFtBCcAHKvFGjLsl/zUBT+xcvW/7MlS1XHX
TX/t+ak45DM7Sx6D3uVc7s4cGs06fqx+sfiQ89iVbhQiZMzY2XzXVUkKRmT5V6eaCbnjsm+wgEZ3
JrZtz1LEhuKc4Qvw8caBMKqEHFY3IwKfsdjTFDRAZFX9IQhfgbhQlGkweLELOrsunp6Pi3ZF9bE7
lbyVsMFvXlB+nudkl68tipniYquE9vT4bldNdQBlFTpAAeYbNwAJ8wcvhg1SHboMsGguuxXt2tPh
ZCvzx1SaKl+GZQbQhnKa5V33cT3+9L6nRMZe39UmV4JgdQuMfJivmdsueFfPIneA223GeUTy2wgS
4WOC8s5oDqeaDU1lIxK1sTLgnQORbLPs4ISGL6v7ElMyrdzYUlQ5K5MasbIyVcEaS8GS1TXJ1skg
R5ej4GzH/8iBYFVxjp8USTtazF00ZsFftHYv5SEImJGAwxuuy87lx4SNW/JI6Tky1uUh087H+Y2q
3kGoVfXI9iF9p1wqOKth0MN5d230i4Eb9fUgwNG98uDi2pLez8n0pYf2CfFq/AbjTdp/cGLaNzTC
7tui3juQTz7qtVFk8f+hM8SiaJcacR1l1rHiC6I/gnvScSakGtE8FUhA+eUyHz/eksNOkzpJRkCa
tWhObXfyM1G34w+uahAq/k379htsoGp59HqjxYkkweXAC5w7VUbwzuUWcGxdHZhvUyMFBkVzV+Hq
4sbSrWrcKMj+69IjkyEhWsgP5IMCmHb/yYfYpbN9NgOuVbMk0QBz0kThkD1HXMC/bbv2GyOeoeaT
9zEIPj4huMQe5T8f8iUn066RAnzMOYhte8c8HAwLIm4TUSjRL8bgzIGQ8t7VuUA6l08OxRz9aqmP
K3A/C5wCRrXRCqTHDZLufJb/V+h3Ntv1AzvupxHRKYAySMC7Wvwd2im9031oSG5J1DXqAKs3Bzlz
228Vwc/Ay/bF8fntpBpTaMH4mYAowTz8XDo1MyZzyz1oC/2CZMXDgxM9/LmFiwU9K8NTndYSflLO
7BqiMAHXDXThyhJPMXMFVojlWIebaEI8Ea0na2numbsNFrrUlEBBvPlAjGfRxNejdWhhj4NmaExT
HwALFdChsZV7jVd9rbkVMoN29Ug9/dwvG0287ggits2E7397cPOQxLGMIF5D/gXKllGga0oiftpr
BcTvkSJU7/epluCtEFaHIMqedAIl5x3mhhCo99eR4MnuXZ9JvfWMsOOGW/05Px5GorNXMJ13ZmX1
8o2RGbAvd6zeufNzvmd9rr+7i+q1rrhvPchpkn/+6vmUo0cTduFJYMOG4rZw49v4oGSUbob9zgIq
zKFyiAcW8Ds9Bh64LobDcuOmw4NeszUEdcjM3DUyYJeGbKbhoToFYwlm2eKc1hAnqrrnwAHlRS5X
lXRvWDn3bi5akvD5C+Q37uPNovWbzt+/q4BwPmFii5X75epwu9df09HMeqen63ptHoKcXiMGvxHK
fI1As7TemWJsSuBN+Ci5CuddTrRus2mSq21f9mGmcmD+t/tFwGj6r5hgzQyEqFHt9dMPDOPRmo31
RJWRVfJif9XsojcFdJhH431xeE0FltYKWS8Ipy4EJ9mX/1GdynLClJh6sby4kfUCdP+5oW7Td6Mz
CBA6MHirdLyBFDHiEZbQdM5G4u4u2/aXbb+oH7z9Ohxz5i624FSTgV37077pgduTxF0230iww47f
IBCGUrw+kSgKHHUa+1WaETxP/BlnbxsARhznSUPBEY09Shj8WVF68Uq18wX9T+1qc84zuDMqKHgl
BiOwL1sYMSUH+F5sg0F9tK8nNTQRgYai/GkEzfpevlfru+lMrEfv5ko7oBn8hmSp92UIqevAYd8E
DC5TFAa+x51N1l/RcQbgH67RCsgjDB/U2grGbmHO0JoJAKXLpaWn/e8m+4ef54Go3SzPohz7GGKE
ho9uhCo4oaEK3euV0djoBe9bznOxMPLGO5hmwWsaBX/vP55ehdQ13n8ZfOdQpJ9rIQarWTvhUMfF
vapezCHjpcYbRkacsFypDl16OCJx2bYkPLDtOzjWHEAcwEswCDtXkQobV/urL4AWDTrZkksHnr17
XjzXYkxPhjhGdk+DY53p2KGXVpMwhzm3/MW/tCBtidaUi9jC2qnb+W4UEaSK7hIZo6vub6neb5q8
XNHJZPLVDHvrCJ+m+l8A1uUJz7YHc3WJavet/A6jmUI4TIv6p/LgmbYChIW8uS/9S+7VZOH29gzB
thU8k9hAsEGBKGnK3PYFzEkPADpeDB6hiSgu/qsp6v6jgK7ClKywy03grARQtm/l0G5nHGWiP8xH
ujT8zThO9f2degJW2mrdNDvlT8nQQ35amS6wHT5/6XTJX6DntPP91imTjsUga3bNmWsuisXW/A91
Xr+dUOm6p6bjJ/cxrK945+At0O/jyoXpSZV4zOXh3wc42OR+CAMVBLuU2po+ak9h/l4YELXoVQ8v
sSG1D+VZrKbLsR0pp418W2O8xzdSEaLNA3u+UtKh9cQ2EhrV/+hgscqjYmAlM+sJv6gF/Vt6Idzf
OBF99aUvNULSTv+9z472Gg8cKtJuwJ0720XEX3KEMQYz8v5Sojos3Yli+9OoOZdKct5LQl8u67gz
71ab57/Z5o20tla60pIydgtmYKNEMgXz5AewPHAzmSweoXyQ58vmAwlIZRmmoWp0Ue1eAY20ZLL1
uOHfD9ELEyWpKgRzn5dcm342byoe/H1xEmLrqOK1V5IrTf9qzCxkFbo1VLZlBHX8NRpnHCOzKntX
/PxGWk0lfbqpulgkVsxdXTTBAgMKufBEV2KM/79lbi/wgCPtdEaT3PoL9KJneaON1NPHXsU1vmPg
3MCLdsIeUOLR7VazkYJUSPycQOJFUZrb5LJy2mEYv5tdYhes9jucZfclLhYcuBqbRPNOqcKIw5AQ
CNSS2ubh2IYbZj1iVuJ4343UoVOl+DIaAju3ngjBn0M5dI/w0nXuNh90vUWpj2emO8p8/lThMATl
Pd+4Sq5MD+KE5o+DTVze8bCY0tnWwa+iG+1mH4tx9mnZyNElGv7jYfg9qu5qAYrzpvhocUUre/po
wN2FQ99DTDE9VIWcEAhalrZBdR2SSVHIjn38mai5XP3qM2NC3pX9TGQwPt97UVaDXcH9mUfcvJ+1
aCJP84wc/cm2/LFm6eZiJnOXAXTF/GE3KAaTzI6iq+1XII2jktpQcXkUHTecsvHxxZWXLqrMPHuI
qv/EMKnSi0PozHx43Ck8RAsbBa+/lkk1CNLlSEO8PyD7Vt7IKfX3Ewn0vaIA3x859muocS0yI/Kw
GWkC09n8Pi8HNUqNMnlZWj3Eda/DrG68Q8ftIAwx2lWGTfyv7+oPS3SIyJbGRLad96uwHTG28zAT
pfiiWhvetd3CSGLIFU6Rqjsug7UmssXx+BPjt8ygB/KaipGwbHrsGxOVKlnoRADgN8oG6wutpUBa
jNf1c1k9GeEIQySASjUjDSDn5V5xMqiJz9/QajFGnmuMwBoMdciBIMSWCPmLphX1ZwzxlPVianEk
Hkj9U0kq30xCGj31Vs0iGZD0ykqZDi+kSi7J3FPyQOm1dJ6aYh+Abv0ujzRveYxR7yWvvXPpvx4l
ucO5ZtvTI4i1zYBXnP4bVwnu1/2c4kbcILY0k3l6wvP0aOE6YyIrB0YyNBCG9Thok1a5b2v7AsiR
PHSnRxf6YQ84tZ5w8ZKxMjqABtZeJNuhqUxkkcni2EUiJu3TJirx1YjDxMCjtokfbuNZQLyTFCMa
wJjGIEVuzzVRmrZaHKlU2gA77PIHsHMGvFtuZ4xaDfL+ITTNMt6LkffJgMyhPmBVfgZx7mD/Qjjo
nwlrCSBEE3LhLhwunSs90sIIK4S7TFXMD1tph346kfooxDOVvfw2Rj/BZYYoWTeqRoYbv4z8olM8
xHjEcS1CUf7pOhCm9bue+bu0Huo7KCHL2m9WmGtwpUUy2TYMV3t4VVsa1VY4qGbAbR0UsWbBTKl3
A9g1wB3+xr7tt99b7BIKihMRXATzuXbzYCExa8Aa6eihZVz4tvyi6iOM61mmsrNy9RzIKVpFX9bX
PLfe0qA9klw+cIx4unBj7mxK89G982d65OSDSL0nXHimQZgMC5M/3qVsilnAJ1+DGUczmIIOALSp
uvJcAGjTJug1JLhlD6aRa7j6b889eDG2F7e3m6DGc1zgCcs5DAhqqlgWcD6cudYHy1XikGJ1XEKc
i9C9Lybe1ylAKJQr4sObQHSppK8yJN5YW1R3mXAAiOOXz292v3wqK+txdi2oChAvr2ey41vjAC0D
l6KTlnrhBAOsnbmmBgUltFNilJSECTzZfNSwSeLqDkvLWz9UL2SIUe6dw7JN6rswKMb6T4WkHJpJ
bM6aGUKJZ1ARjqi/ZIJCMRW5wFpwmmxJG/meHuu0trbtULxUpWSIAQJA3TWGQ2Y/wRXUMgi/eS0s
BU0kdgGZFWW+Dpy0UZrvumgOugqx/WMGiMPRaUEWzWjqXTnsdjjFn3SRakIrDvBaepDMspConPG9
FjTzauKokt88v7irdZiWnIAsRbKxe2MA5TZXb4tiwkYcioCM5zkZJ7cADdi1Gtlgcnfw6UGlwxE3
Qp2RXJE4KQw0klVmMHNm1rXymFnhGCJg9IhFfFjGRg9epdpdtY22MuQr5hgHUATllNtYK+M2LZG0
2UkpCXmFME+htgGalG3SI2rcxzL9eQPN8CQUsryPzP9f6e0B2KrddnTo7rzvA8AdRim5ucgXNmJB
qhugUHnc7LSyKqnAY4Pagb45iPI/+3r6Dm3BKgeF0MpZnKczW4UWAauoyoy/2y7BzbXwzWhPViyT
Z8tz+9vNfCmzfxqJEk1cptTcUsobUZ6JTVNQSgLIyoOsqQikr45Ccbpem/CdeXwxfSL8JnlHSrPL
wgCC2j6hvkCcXFrT/kgSEjf8arpsxS3rY2m675OLnMPEn03tWUFLpj+LPTlaLPxZoE3V92dRDLcg
DaQ5yy2XuGXZjS4wPYRJ1dm9lytW6loyxJqMDuTBUXIoi8lszz4QsfC3/x+0idOsjUAbO6bccW+/
Yk0zr0By46zsq0pRbDmYBBiFlubQUmUigmIvEudQhQrezyqs2FFikowzBjYCxQ6KV2kWXZhUr9UV
G+sej9pRiJB3vYv27b7vVcCLdqpro+O3OyWJVthYaTPjBbRiaqXAMliS7DBgbaWRR0dxmjb/62an
49HeVaQpZvrShf82h97AECSj9E0g2BRZpkr+XszjaVe3dHItywygErxtEi8V/2e4J28VfwGkiP8b
+xp0gjrCFUTLt2itxAVe3Vkpkb3g1Eo92ypGcxijddKmRdE/Bxk3VEMSHbDq3nqzm0ijWeF+ZB9x
dt+zLzuHX5RtM8Q+97DOVIyJVZj0ejjM5CKYAqmloDS7Id6OTWgr8m7fC/J5lZGqZTa6rGdcGQru
5nIygVTm4DwUY+vvS574hF9RjOZRLfoa6uUUdubOnUBqAfs3db+UjbD/a1vJc7dKfUkjlQmJge28
iHOYgLo78jmbUEiZiSJsPwNOg1muMGAjwC+F0S0p6SpnTFjahneegXMqrpcARSBAmheUEbKwUCx5
lEkW0KsA6DKPRcmhZEbhhsanPDkvpm+/3eefn7LrAhPbo82+zOfvkHzNFgWKgBfzZPZowXmzTTzi
fkkHjEmmrwzaVBeeCvxdMh3iqYG3xJdTznxqYzFGHM8Nk+A9tHdpa4AfTzJB/Nz6HvTQapsZiBsW
dwPTJ9VNg0vuIF2n1Bz2i5xbfOPUQ+eCrSsku6IOWPTzM1e3bIn9L5Nmv/ntutZEi18+uKFOxnel
ezeJlfCDeSb2AP2sogHdWwT1kGx2SUSNNO1NtaTbwPb760W9HN+NrbXy89wtVUbNXNDN+3Pfl/Ge
tyfJSyEEVG4QXlqp5kZ/5stVX/h0K9BTVpKjiB5GarF+OJJb4zeT4DA0N7Bx26dnbUyfvrCKn5rl
wl9qjFLZZWQKUuvVgjMZql1iFIorKutjqSkuTuSTa+w+1S5AuFqDt2rJO1S7JBj+swiqGwmifA+X
DWCIdpBKvdA6RYhDhpGGIx4A7oQspR1V5+SwwQsMjiWe4YEeLU3SWW2RMDZPW9wF/wa2Rv/T4y3v
vsbpKbmse2zcHteL4I7GKexXjRDeZNXwR3ewNzwUpTfGReR7fGwhi7UuT0riEktPeM6ZN1J8CBtA
H4V1nrzwOP1GO4NsBTSyyAYN9nZcADEQhjGgKjKsHoW6I298EurBpKF9sfPnm3Ga0d8GpDSi818J
U0mnoQXegVpMz+wqrdy32UClGU/BPMJkoRfnrEsFJaaxN1TIskw5mAAXe4XnK0lxL2u574dmSeN+
aY2Z88X17XijNQA/rgB+sjLb/Z0Ypl2LLSOu81GJkcoeqnCYVPAiz9aaXaRa1VEyUd71jdz7VkDA
tU96+28dZ6CMSpBM2TKnCBG7KdWOy63mcDOhGwqvrwkTzur2YBa8uOdfTUIUBHFK1kI1MjA35GlD
lwZ8jk9zMtIb2hTWEDL7yQ8b8kMNCDANOheqo89aQjiSrvuSReFwOc04q0afgjEFJvTw18ScIc1E
xWJmZzN+gxhN0iBTczX4YoCqgJXFEMVAt6jBWAd/GvSdKKQWvMotdZamX/hS7XQ6ybyVEkLeAOSe
HEeHd/zmUOk/x65tfP1ZCg13aBPHFn3BakBMmcAhkCU+ZV+tcaFK2HOkRkkz8YuX8FCddwRtPc6d
vS08s26KkQTdPOZEgh7frMueZTfVclSBryDxSolUQZBNpDBwwGxLOIppjy+cpuql71HYCprE5mX1
iWwK01/4LGxz1Mt8xDHzjqMt2AgddXeh88vEoIQ0Xev9nFhbrBf0NjlPPNs9/i2qCQamILsx+hWa
7UktlOxxKYy7PfGKGNhnNEh527PAP7m+pIuQy/MQahRIlYZ4inD+kLbIb/w9RLN01N/A5vcKVSCQ
FtKhFjjSKsyAKiOFz9Nq+24w7O+3ASykivB19ODp615V+S7ZIJIbDWqVNKaUefJHhUg1HI0kE9yr
FutWLvFvmvM+pLPWJIUGLnxs2HzKLUOjdvRdpJ2zAazZU7DxdkHtOivI2TNylSoR7XFboTcWdDE6
QMTPeyQ+gTl2WgJWg/szR5gHsL/yPDDS5av8MV6TroAuEL0b9ifnncz/hi0nBYAvlfg7nvS4QCTI
0NXcrB2Y+rbNyb++7du0DVN57eynd8sNLHGnY4WNLhmUVFv5FWYGaTDxBPVE9IREMNsCbAB5dCO6
ell1ydva50YvVZAGX9r7qVbUxvQTzavouS8OzqumPw79kEXltW5lWapof+nrFNkQj4pNp7v3CMK9
2GhxCzApf+9oV3uxSB4dPk+s27Bb8X1BRKoTGBFfdJlowUUfnxgyfyAIoY3hPN826c5H29EPkaIL
BGt/B+C3GwdQ41Qw/VAKfjKB4awO/WlPgDepd+pyT/WCT3v9pIWvQN3svpCNR9oX1+ejAOlBlcuH
VYvnPiBHNfcM3Ul+nmXHlvrGNzLmsKDDOGYy5ROl2SodxvuqJ8NkoKwRCYjihi5IuzSx+frk9X8e
T8c9+3vV5Qdds1wgLvgc55uxb2Stz9iNnhw7eKFZucsa+U0e9hFkcmlRR7zDaB9XGBO0lM8yQm5g
C9b7gH4Tey2gPRlfXm8RgQMopb8ETfrFzdbEnzmcSZKWZI2BV7n1kdAa9qOe8ohTlr8BE5Dcs3CE
iwV0oPCzjC8M/uQPhFCrCqwlnU3X/6v1eEo6cExB0hdUQT2H1uHBmBHmH9sFd6IweRO//ECN2R+M
mCP+s4aWR/+G9I1GvWd+khagZ6ZsImL9MsaYchGXuQ9jJzz2Hb5F8fFaPJ0PiiI86wxbuXqkM3zp
mVC1zpOaJwg4Qpx9Q4+WjYFakxpECa3cvCL0JysdB2DS5mBVwcyBeLexBA78121RKIE2idGRUrEe
LVlNUF+WKhtIP5YE7pyjHzWTfG+cVaFDet1HAv64b/xzrsgajbjzWp3FB9fhWnTCR6tc9qIfrnQ3
zDjul0Op+i9nKpuTjcBrZMd+ipC1ZmX0LbH68f8WIflBJoYWK7k/GNKVs7HcCfwaZA/jpIfgmEJT
RIIc606r0R+dMqmymuUaqfQb1SOWPy9Ish1Tk/c/rX84CQDDWIE/X2YQJCUve0XOWE69FC3p885E
QYIwehq/eAprJz1HZ6PiRdsqJxpamw8yADQcxWuFKOBMdKHHHa+3Os3Lo1r6P5QZHffUhBGRQCB2
TEVM9L17F9nxRJMoB0ke4sGvlcrPcweu0/lxAtvq3EscvBrfGZXWQ95ThM+CZQWYKXVnuYOrAFf6
mQYCJEfRo5a+kphf5zT7EPWe9so39R0dt/b941Vn387SCQnLOBE5BfwdT2FzQ7Qhf7P89U0RR4Tk
N9Le31o6zav3PjeKgHO0qA1OKQwfYqFpBTKMexAzPwoVxd699zuKqDbCgd2V/aB7KvtSKL6Bp4bX
R4E6d6ISxFnFm95xGvTRulaad1sgx3ez0ZeO8RvWchduG6RlMIoMdI5Vjzlj6kOGNCXhfzGJlUk6
cMzxqiUPIsJYmvmy8y4IYz6L7LVs49tBmh3clG+ERSoB2f00tWtJkGIswMs/epCaPv5M+LTcOgbT
YfqY9/ClNb666eYi1ZPXLRO2XVjKp8MqROiDdzDTBD1BGsBlLjDlx5+zh0FLUsPs8YBliQ71MjOz
IHTGPLFtmGYnXJOQtug+HApRQF/63YsM2AP2vyNt3qQ4giocksSJkMjuHLRSnDRbCTnT0UrCbiR2
iqHyPpjVJEaeRk8gkqdgtz9CkEpkn20DV5jkcEMvhXXkq6N3VSNYlY2sPxzJ1M9CwKY3ISXbudlb
2QX9KgMDc1sjclfDdxw9gdRW4/Yrym97nd2Z7L+Z54OVrcU4O246/BKOVJ4eUekyYgiKKK+yxgYd
pC85/SnaHGUPPDucESuLKe8bsF473neCIqQiVf9SAx/zzHiM0UcNjeq73UfsA3nB85ZWx8bsbrnH
W1P0aZGyqqMDyowKNqJITM7FLhg7yAsMq1o1rTomLRpN8UAKWJamEQE3uaKnc9gLpBReYGmHqHWv
g8mPbqpXQkXdZv13EUz+B3Fq9m7AjhMj0XaK5XHG8LM0Knm2UcfecMbBES6nMz/VmFMkWCxnZEUE
MXU629DCIB2Bc//b+XD2d2aLiwEm/MAOHjEa4NbLGzyGV7jgDIFoYoeMiOCw+U12lbPg4/PnNaix
HxE9FIMhWONEwLYrGeaV6Hwnt7pLs/rbRcn6ykW4Rjt1BqQX313wjOetubbEmCkzsW/OeiCq9pfm
XDKKG8OW7dLI8mOMZN5kOoZcDEPcAtBE4kJ6QA2Oz9UqGo2QuVT5m1BvLvd+8RS9gnvvOSVMRu9e
n+hipvUEEWOqS2GTF2I6sLYIGDqUiurKMAg94ok7iGfVnXy1QQHXjr1CMWowYCREiQzXtZ4CW+Ka
unIYNfDuG6LjAS7nzxDgM/ccw2DLSfrKr/TWSk364rh8D/ykAqOEeZqfRR4GZsnfT3aMEmmwbZCV
8PINSx3mcePKbU53WRgHZkyeEMMNHnIJxmYpRRjLXIX+VWKTDo/jD09JxjBDVQX6K8w2RlCaTqny
4yjyiR10b5baS0670TmASJ/39WWcOFJBXMGUPs/QsLcFrT1JXeP5NBcDG10+ccN/9Z1mC+Fo/zJD
h/WUW1ZYHNG3XULH8Uu8jBEq1uHisFnwv2St6x3MvV5RCy0R3r9Hd4vVcv0CRKj1mG6+pcvWyjJX
KzoIfRd5JWfwf834MEnJtmeWOdB5Ly8wGMTNdo8UdgtoHHBzVjdXIFavHonV98ai7KC4YVeLv3Lh
zL8nDSYYlqwWhEI+shAWyaccDRSaa8S41+M6OqQDDcKxLrF6WVw6atLaGnzss33iB/1HKSZTl7E7
LmbzppvS/cdYNaE+8yu72y3mQccZD5vp+kAdBDopQceetUNUxaJAEItkwipBbB7l+v2+0dgrwcaf
ibSMO1okZC9L9L92i0jE24jZskJAXkY617DApyyW7w17LwvhiV4TdpaggmLDOn4c94Ac/ogEDcv6
AKaUXxIlfDfTOi5+C3bB0uPjuX/N9J5Y55ERlwZ86K3uyuzNBySq93lxsYwYAC9ap+bN4s4GyyfT
Vs+pQd1I6EixoXWwZ5A0W5vzmYPPTlaB1jwvhDO8zvrcDZNS2+QZjNPcT/zwtVn8NESTcEfD4pw4
31hRNm3NE7THjAKRlXGz0dMMtlcxACJ+71aXFCDfM/UQTftZQfq4d9HxRvUftVumWp5+sQwZkd+9
ceGzvypnYlxUHOjZbsTSdxuTSZfo4XMiK7F6anwoPfn056z03FfgKSpFr2zBp5PPHfRVdKYaL+Pz
MWNZnUfCTShxi/QMGy3nZP4PBkiMpZcIm2GzHdG3e9YTorGew3bzJjmPRc5RwRX39IqTNl9ll4KD
1H31t6Xebl4fm81epkZsT266bsEdzOgL+X0zEAVBtEA5BavD1kpsaYEmjV8lJDTxMcnkzEieDd9T
ExEiioym/6joASyhSQ0Gnl6sTNupYEs/xp5YWfmm8RgjkxBBNJZ4JCwmD3YglnR8SFUNZlh9gZd/
hONnWocccLq5qRvirJSs7tWGsF6y3AAJ8P/Xcv0Ex/p4QJfqLCeGIzXrGyvHhBvGK1bd+wVn/EWM
smO0sojUK8M2VB9dHkgKagg93spNdx65HtGKnFwHnipMdgo7FgrYQAWOXt9Ws1rlh9uFAWKXh5s+
WdAkMXHlE9Px/ps6PXAgOgbihWxySVfks5LYdJ5OozPPZ9k5LR0daRE5UHLWbFBMHT+nyd3U0BB/
+Ou/u7bb0VX7yxSNJJG8GvnKRpZXLeWF8hxlxcQnM9aIJMQVMStDmjxoKNfN9/X2oFEBFJ/wk4LJ
QP5p3ShOJ7EYACYnKha3mzmYiRNHGPovqwcU19lhdNoKduttgTXjbMeakq0dP+KlJqKomGb8TNAz
ukEaMQL6ClQU4/RMhDV2DnqNZtb1pp2FmQtc1ZDLjWA3a3U0M3sKutvd2EjHXtzJnJnSspRqx4DG
YgpRsqtrbUcv1vmXVlkW5r44I5hyGrMUbZB+imHekIdOYsjQSak/Ecz82SmAHUNizX1wrynU3m7m
rdILCa1eV4IsB1Y+xy/gByLozEz6Ik3k3Oag0TgQuJsKHYEiGl3CBZBuPS5WBSQhXb5V+G8KHS7B
3BsvOui/kuMSwQBkNRHklDiStoFpSk20P4M8TotZR0eXMntXZbghHnzg/xCYLiVnmEKZcAyqE6mb
HMwveA/VXicYQ5JniV/1ZD3+JO73IVaDy9SWHNBdH3vmpzoR5BD1+YzYhOLSULsWMDJo91v4QW4D
3oclBtqGSjHr7Hl024iocwkcGplNSHts7nRkP5qN0gyPI0nSJddSOwzPlFi+Zqbp+ny9/eMtClZG
o9F+DRgN15NJ6WrWGnguNtc/LpYfov7iIkC64XiZ40uYpPA7eZcubKKTCP0nSrirlX70mX7rA5cV
eAw3t3AN94CHlZz+bSb/nEesBaMKXpRn5JMqK25v/dsAFmbufoWgKvzt5t5Q20JKkeX6zunMYKv1
7Z1S/Oc0+ZgdjpsEYAFxo++2kXHrTxWFTlvGzK5uDbqm+lLsH17FJKm1DnXLNxT6Nkj577k09UpY
Xj/9WA6w4y7Jr3cLphH7/IaNrW1Y0JdW0bV8DJOsLEZWgoy2VDHED2z826+Eoe8UQ05CBGTv53+n
gwLsudSdLkdXTcz4jpdUVQOiP04OEoCtpuLl7jq25489z+HVQTikvzY6kfxR3evNqPQJ9spfbTv4
6KEzP0N61qg/THMeLuthi1R4+8CBC+tq/ObJiNfCobZQ81ANjLF6dSXYXk+TkpfS/rd2YBZuT4Tk
SxqxKIgRgAH7QxgZFi/Uz7r01iy3CmJjeeKVee13Gnly3ErQ8Ns8P1JvEwxR3f9EtxSn5bD2CmVR
xewZqgmPymuwS4I8MoPUKQIsqGTw02DkYMDGbAEW68j+2CXX06zY3SgsFvV6B59qc9XIiwmzYdWZ
/3Ur4huTjczIRWWTGzUaOh4eIDpf8vzMrtGSMp6NOsc02EftDfq8toKMbcXbEWkbLm/TyoQdqLNb
tRsBiFeQxTSC5B2NcJEOIhU/fFLGZW3XBamNAtohSHstzEIQf13AycaItKHYuwJrd3G8wa3kBb0j
yDc0GKRrJCeDxbxePimGj+4uqXd72J3u0Zf+3S4ARALz341HjyN0mHTOCYE2fWBJXEI0lmCf6EbS
wdy9jtOIBVjejtooRSQw9xcxRdLQcotCBCA62tGkA9zj7aU8vDg9DcUURAxhXv2OyZMWZ7Z8GpPS
CmZJKAsIbfTkPlq70gL+8GXydOCZ3QDabieXW9+GvWn0bO/DMJYGO21HusL7oWDpjiTDl5AtLuU5
5pgah1jyWxo2nYJy5CEppyqrKCo466+SrR81krzX18I/Qa1AyeJ488L7nSwaNzJoEKeBkxXbbDap
4OnJA1rBlk/y+lcL5ma/nn21xy0YNXwJZYlchtnZEmW/eLt/BQ9r9uK3pkIz9zsePGnwGf7fgg+P
ITkK5f4JR27O3j1AeCxIjY9AMgeFE9+blcqis6jSghSjj8KFm9EZalBg7w8iaYfhkBpEPnQdJ+tX
LZev/SQHYf2dmpCo73B9RxjHs7I5uKs82xMFgBhQSlkZMKP5DLeVbnACUe9ZdSN49feIw+FRK3sr
aDF/Dh5qWEfh5d2RTKK4b3qfqwCo0MU255XmdLe7j7fDnUngxsCJSDTHV+jneU1vw+ZCQ7/QkfPs
RG5YRp4wf5rzVaKucLwVAabSKvlayuWBcnnf0X7ILK6ucnfSu87X0FoHuk6rz6jvgMJWpiqxF2ix
TcWH6TLlbyMAK5UyW71l307gQTyHsEnmd4YrEN46xXqRgRle8ZWX7zYNeVGB9L6vaqUq0dHXRlRe
dDfjVIWxQ2NE13wJV3UZY41ZW58nNczs1EYXjHI+5p1L5VIdFJsA4i+G8RcOHrSU3sp9seKgolsg
AiwX2v4r+lfUV1pywmRnAPd4z/fFvWt8/bHSVLWWvaBINHntkxyFqOx/nQw+HSL9a0vt/v0CSDiA
OwmlFGdj38mnZr7weqa2Q1OMaLAx3OjW2I6ic2wAjMkTOUDRCCy/vuA2r6d6/SXpTdE5V+BAnU6L
GKLQwWGasDxGbBjtyd80rIC5JRSXgj/Vf3LEML+XKzg0uSEbOKcIekzCNo63foRaDmhjR/7PwwmH
uVLPl5fV/x1BZ2FyanODc8M769fGysTdHzJWrcMCn7IBY0bMwTI2Ypjnwg+AjnOE3WAYLsE/E+ML
tCGyrysYe3rzLN1M6dpZHANEEpXOd+/cq5aMgf2cI64JyCC8hNYnU7POLTitDa8+U3I3TPYHwTWv
IzE6mF4f83avE6Fkc+R4JN4wLQhzIRamixCnOfK+8yAMfajaKNsTi5WM1aAhywedcUyYqmzRUQel
7YUEDv4sSmmu3qZbFuvvJEtdG2YleCvlWRACPhp5+D9SINlG+ljo8ecJEjgEhBN2AmwL2rksEMsB
gpb+1ATyldAbJL1TwlB9Jtdm7sO/Z7jnqmehXi8MD/Nkdj1UMILRJILh9YS/+H4f1tvyZK+B4nSV
PzPkffYMrn5Pi6IU8TaFq2BynxaK5XA4vFXO8GrdWH1HXlFDNKLBO+ftNTdKVCdfKEfFBljLbCgB
uY5zXUbjcPa4UX2krv0NpH1AftSRi4Q/XFDemG97DyS79dnvKTRA6qOXGKMMhP7CpMQYnK38LxKB
9JN1NJ4WduiDUdWqMC9JHRqK7BhoPi2p/DBzxH5lkOQcDt1UN/1bQeogAMeTpw/GCKTC57qiCYQN
qTOGEzRleMZunnNFCL1s3yL+DKVWjVa2AlkYcoyUMDI6UsqPJtGa3dbYQntsk9WOpfK3NnxQVTkl
Cc6jKG1Drelj6r+3rhnEhUwQwIeMmdhEiZcmBk92pvb+aWuH9Iiy4z5J2xl/E11KxXjKZq+VXCBi
0+c7g+AU0lTvkUxfCqNFjUO0IJqsUjs8pbdFch238/dBtA7e8MviMpjENcQ8tyq/CDdUiYLUwdTX
wvaEFzuUD8z7zwTthmd1HfOoJtrwxk8reXSRPkkGTxFFlShNpB0st4/N4TIwFRzBK6JvHwu/xSat
FJdRxwoqINleEUyEEOVyWaUCJk5rp3nb3Gc5ibMZjK92D3aSKZSi0B8D7Hic3t2dkdOKWfImhddm
/Di7UvIuyJXgH4NFAlRC7J9Xp9B4wF/MqQAZyrxQsmGzDHWwse2UvIuhTMjenwzRLsX6qwZcPp6w
bdkGTdZ1hOJhEUzfH6BegY7NKflVmJ8im4qE2eXsWqyc3vixjOLJ3lRtRDIuCSSBP8eDZe/f6JX/
+xVPfJCd0hFR0FrOWW2INfFn/jyzCk2wHwYtTc28P70zh0cNKxxe0GXE4FZRyHDrXd/c51QJSApd
R/qsoncoLR35ap9G7Nm7fCrw9aSlEAr2DySxWGocr9ma1/wk33pJIZSiZxFV4sfbX/h+toT56ZaU
L96u4ik1zavbyWBQsQproCL8jrXiqrx5/bhM2xVbJgL+mV4FMhN/POKZ029jj3+bcDoXrsFjEczo
yCN4zuEm5zbZnXF+GxqekzeZH1MvWoLg7DQRy3rNCOjBw7sCPmfNgnQNVp1OoeNZT75vojh3lEmu
8wsrFTjVojgh4Mw82sVyzre+IGszw42k4QPvkQZ1bfE0IPJJwQHUOQY3Xdk2ddTsQcUhOrqFVMYr
IwEzx7GyFf46lVi8TvHyv9QVHBUTpvVKgEPzgkxjbP4KAMbdDAmUWqnbMcV22brsdi4SKkMe2HC5
+PuFVvyokG+4e3AiudRZIIYtE9tlBrtPxDtnX0MbPz/MkeymUjd6/xQ0VkkhNP5HlzPYu6ZI0Ndk
PDlyEuFCGEyZSCQ1NCwSSTsMdIWN5HzCFJ24fvyQC93mac197MRnR97wmChj3BAyxIwWefFxF/zr
EK3HFcUo/ewJ8RLH2aNkmHHNtLyNfcMhBKO2DJrzMEsCf5TqDx2Em1zzy8p49Mep4m2gt+Q3NjCn
ViRzEcKtS1INiJJTWy2iS/gE79kpJu6pLLXXdgxs6dPHEcl5VnB+w1RTz/lKnM3RwoOuVPxkbZis
vn5skCTHfMsnEdz9OO7LXtqWbTgVDOoUCfmURmVHE7BUjCzflr+geekPbM/92D9Nf3194SyZusmp
RR//ojXrPWbtvEetcIltiYFhcqIUo1SyPj+pwSAJA6Dsm/OMlxVKXTl1SzY5MnH1XArFHN75+msM
dISi6lsDQO8kFWp7+SIvA9QPAxpdIEngqUXHmbJ+D0ZooIl73l4WnGYc0hgRDjRwd8IH1cdKSt6J
AkE19JEDGrDjUG0ot3z3RXIyEYnwgGJkN2ztTTJx38Hr6dNK+DqtibkgVi5TF7KSBuzaXL2IcV58
mkQagbf5iSPl+VHwx5YPeqE550oOe/o3iWPxBOZXw+8V1G+g/+BPNLMtMgSVsXSx4kn98eAFv8oE
SA4bKCvlXo0gMFggOydDRKcQ7JjdhNHbXmTMubpOd6GDU1NDncTQwbPp7lu6tKwDJapKgOSO2daQ
BeHPMxaT9HMBkxZYZXZv6nisezOMR1v10sGRIK1YSw/LTGySyw3OT5CGdJ4QM1WQ8okJiPvd51Cv
R+U7R3EJYyzjh66D9+tkBlW0hosWNXMJZ4bmWZjYLAidjFws6kOnRmzvt12+tjmG5/Yg0RZvdkWK
umNfE3ghvOqi/ZQ9txVFLQZMl/Rc+jaHXVlTSbyoLEduOyvXu8g6m0f42x+/pijkE0ND+vCUi/Dd
MFmajPEvhMTq4AsfR2B9fQhysc5WUhjQywqlygHl2N1Amzzg7Pkv2Q1gC4A5ovYBWLo8aMeNMoKl
XuX7Ms4GVQ/x/o6z3FrwyrDGx1AewWUFFY20JTd43vTarT44CPlGsZ/aAkTfcyj/vCe8Q+d8OmrL
QQauGvzjTJKLPgGuZC7rrqIHQ1dT6TvT/xKdjigAxh/NwsJJkJcVtD2idtxik9Pkc0AZhIthmCp8
FBMk59pBelrIqTz/hZzeCJ9Zf5Zbxx3zz19mb97Rb04v2EmX1l9IAvnY8JcYM9sJGXBC1oNG9vYq
V1JJs4+D/kANxJOa0RxVuxtkG0WjJG3OD2m4azgFdJ32CGqUZAv0dzCbWHGR66UdqOE/w/jBCg9B
cCsoqaCg7jkEINNMk0QuM1xl8A7uUbrmWQ+rT+BNfsqppWorCbMf84thYwJB8aOkD4BuRNTbvhzi
Kredtg9+0yf3xHdy/wLFPP2xqLxNmhND8ozP/hPwO60IpOkSgbQmBdVr5Q6RRfsmitGVIs6t86qi
UI7JdrCQLGYZDirhCjmdgnCcKdp6LFq76TCG9iExHyF45fBBpMCWPM1uyBXEYn1dgQCMvRwzFm+A
Zd6ITXPguHeFIOp8qfejljnmB+MSrVIVvroUaBhWbrTRnxjVeXonU3ja5v1oXzvxIy6UJ4gYSzTi
zJDCrljBh2a2ltoj9qsMZCg/KS2Fb5/94k5HoJQU6HMjiF1GvpiW7kBmjOhaQk+E5cXS/PUQTcNd
Gtm4+Gklsyj0wwGlgVW3q7lPkb05EpadHSAXc1931rkGM44lqB0IWgVjdQ+h+0kmMsnLBBkI0GA8
NuCbxxQt176gX5GVcW57KaHrJ/XaT6YX81pNqf8jMQJtuEl3x+2ttioHfX1a141F3JmDi8uekjc7
25LQ0U8CLlXwBghOqPRb/K/WpB01vd1gtqzq+Y/8BrmvmdyMCshcayA320Bydt73sINIuxfaqZh8
0qd1MrBVM2V32Btf2l1vMmdiXnAnpIs/mZDfJReUguh3pdO/koUWHlSxAV93p2dx0uDRg0+6FCUu
iW8vjd+02VHuxBaKjPmm5H2YUkwkXA/9K9Riu72VjbO3MFJIOCqvuNNHx5Zoo07dxUNRZUWCaHZ2
Y4JuSotSYDz+ASxxuO5NZ5mglWg/RL9tDo6In5J0jx8cQR3uDBXHUnbkBDSom9QDS17eawxiicYu
6xYH9pC/KCdHNcFp/GWsu5+GH4lT0gsU7iCpJvQ0rMivDzshnaAXfpT1UmKx29x/AijMz1ButdXt
E263XBZb/v8WZV4I4EJMAbyB37UBdtwmMhdwzQC0rLLDraKGo9Sf34EpMJdVpMmtKi6PZ3lhCUSt
//kr9drUPBMrIiclgYzSk/cB48zXDJBwHnhn4RIYzq1Jm19RM+VyEDzj4gt25B4zFZSqWw+sNDnN
mrtdVqu8vPKGxc+AuZSqF51+rIiO3dkGRXv6cnUQTzrcGDz9iy7CL78cAC1cDQeg/+b1IopKklJx
L9UI1xkVlTSowH/2+bLrj+y1ELQIV1nKiBapHxrLHnlOFTRjnJVMvWG3LcQw/H6SlopcEFCAJCwk
W512Ek+JaYTLl1b4FaHIZ7G8MF30zbeyGdjIf53Jj5TuBk9+PhW2j5wNj3Wsh1ZxB5WUyfucn/j1
NeCwFu8uF2hnthTthOmGGcixwnnX4Lk7BC1GxETmG/oUoEfJYN+ZREmyaGhNr9+JfeNdaYL4Qi4x
3uvGXXkmTaNBoYUt0WSijvOeNBbOfk5g9UGMU1+qBtlhjWz7n2MlJeeed5RAhW/5xMOhkcV/aTZx
JRDX2royvHDC6piI0pBl2li0SdNU5PkDETnGqP0OCBtObiJzat56o4hsz0vTwWDarL8hqCkxonjm
CoPFgwkuUk9FjbcQCzOMMLDEBr3rGa9aZ5BbqZvA/sM8WJMEWOsyYBUeBwTjYQUuM5g5WfGldxMc
USo2P3jElFjeFkb2CaU8U/PbcweslayrgDQFbeBvXU5+wAqiBt01unUMZjOIprlRBcnx1rCat7rd
2P09MuNyOITiFrqTf4roITysKNkpD1Htw/GvQblr9zgKr4MOT1coBqzZWdPMcqyhEMxQF2k/U+Eo
ngKvVBDJb1LTCdZL2sCnPwvhqyo9R5NOE4RXMduGsxKkZ9GEOXotM4IRJSf0A4a+TIeS9Oehmeb2
yuUypIrsexxPAm7E/dqHNOCAac+QUcEq0jvzZivc4/spb6XxiAUZAwtujrTzm/Mqq1v68C43IwJ7
ao02lpaUEefjFGG/WejVZJFH9VnStaiRUbKjQputnwzi4ks4GXitax9mme79nkR+x16x2vloGdSv
I25tqWcO42BskORB2BSR2C3vdMyKZ1loEYXa5ApzHS/fS1+iELiK0Zf+qrhbAsBYjSze9qhnqmkY
EVwI5zEj+d1FrC+DH0VDQXcpQodglOo7xhIPjfOaRtdaAUrMbakJ75A1nM102NMmKA6KR84HwOQ+
+VRpuE56bZLUmV0FFdM+OyZZZ5PFkQ/z/rudCquTi+036LGXyVfsl0tJ0d+8i4aavgEt8/N+7xKP
y5m/37SNJs5qF/SjjNzCQE7RqQ+GsV6LNgSwMkGSdTBrRyYZNjRXQfJvQk6faJH8I14m2BfCvooW
OXJR+1BjSPvXlegDEZ+yrp4G1+lXaYIiWqzcVpFTHKR8uViFouEnRJAuF0Tr0U/BqiAmsgfxih1f
GyxJ+ejIOyjqxFqu/KS0zaavM5Te/LsbrcY7Nele09i8lLebyMUCz8zvFeSKmhNShO1fvxNNDNjd
9rNlor0jJy9F41Ykapx7WAQdCC3BKYWJlKUt673/G0pO+Ksa9SgHS/KXdcg0quVlrtWYkvERxMpB
bf0XSd/IzaLjgR0y8aIYXrUsX6mQpeseggP+WhdpIJWCRSoNa76H9lCF+81DhL0BKnDUFe/riZb1
7crX3Q0F6ghWqStShBqv4VNSEUA4dQlEhRfoTJxad8dDBLuTcjeiKrIZBsVdPLUrnqpF4jwoB8Mt
6W1wy4AuLLk0SjyOx+Uc8dvX2p6ewqkZYYBNxpV3BUN+r1Ch7Grs4/RueiauusyPQL4ni1+46thg
eEsfA9eL8D7yg0NzKhkdjC6Jo2qla6LJAVtUjSpcDxDLf3sCsUGU8VGfataePVSQpFygdeI7+aLf
0Y1lirEaKijhDJgWT+ratyDTBuN/71ulOiG0l0UMHdpfYbYyr/wDLrX7FUnhB6uMXUAJVkU/LIJe
rTE69wcvyz6/AbL7RHXKoFLsRx1yrHIpzSvT6K2kUDWlQWF6aG0LaPTmWUmANClDTM9vwLzwfHG9
0SUZPeBz77SnHlBzQ/DEms0xlJJLYj/udGn/23he1IA44S382eTXorMlYc3+2U9bAQvvnnu0e81i
zYUomkfgDl+jwxIAIliqPdiIruDPR9rL4t2DaKWp80YwKzIdVtjujCZsymIZmjczJsKPhqunG108
rtVhMYltKFK3AObNcsispo2t1U8B6019vdsP9nVPj7huF0RJ9mfhkjJh6tMY6/id2Vx7KAMFxBzg
0Mjn7Y1GY9giFEiaNAZ1oMUrkH8AqEID/jzfCsL372gj0/vE6+jM4H3iyh4a1oMHeJ1BmniYldH2
LrMRAN+dbaVnZqzeML4EcMMI8s7X6IhEdwG5GqSg39Zy05INUgx0/A8voK8xJGREMISHdnOQvMbC
qjQFQlai3rOKPNfElyObsXFqBMhWR7HqBmeldLH4Af+i34Zm7Ke39Daz14927XZ3j2tXnITJYqeM
xzSt2Ic9OAM0zDrOeNSwcXffbDwRJE1yJlfAPS8AlqmLzJtr+9NcjMikIVKzmqIGnKyI4L9NGVQt
EwXiyB90CrbyXa4KtbfEwu1Bogx43D+E+gBoF6VBFvGSHAXT//416y0dQRQDPBzPjFXwoR5W9lbL
BhfbXpf6l/Ky5ofoCXOpCEDNGgOhetsNqntDyDH/n14cRr4kSREVCYFD04Yy+O9VnACKk+P5S0tq
sEQj5HqYqdYlG2RHWGsJox+FGN5QnlW7r6IqV/8hI9fRvszEsg4PpS6WFZu7zrWVKzqqEId2AFHE
YiPRFb5pRInRXDR4swMy/bprAtBC+DQAkf1vcyGzG8i7mConMNQZJhNwr9wi+JfKTPzOy+wNXQrv
gf7gIrnfjrA7m9ZTZs0L/AyXAqp8exauFW5O4zrsQcBfJ9unIyhSeGahstHo91276mnkNGKsAnUE
pfatizfxoSur1FyTz0B0xhthfPbjH261qJb1uWnE9eUEFPlVfdVK6isEiGdB8bB2kqICm/eIzQeY
fIADt1z/T8ToaMahIhWNRIi8UpBMzuf92rVG1ggnhtF7mZMMZuCOtTE7KjAxZjGt4gkNmbisuX6W
2J+2dgJVTt4SPOSCV4OoT5X6PJkscdj6bNZ7IQ+K+l9KWAJYgpDmC7K1xzpwXfkZRMRFn5koyq2X
AQO4viXzS4BoIWBvskfmCDLi/bIZw/ZEiq2CEOXlO6hZZV77TxEsWq+me2qQuE+F3kQJ4d4bHIyl
O6atBOp2wn/2DTazL5DbNs0sm/uAHx382BMOCeZJJ2zHVrZmj+HCo2PIa5/mng8JOUGJ5AnJdGD4
+TY5RYXgsL30hMZ0kMuzc/meyN+QjcyhKcee+xdbnoO3Jz9JVYqChoYL55nPaAMT2ReYRaMrS6Qc
z9fzap1+UwLy6YGuqMkYAjkN/WRFW+KWQ9OLLQAua0R1ZNO6yq+QiZSRyeWUQ4n4S3tpujhFDQGq
HeXCV4N9vCwnSBabA/j98yySr42s0qAOgMlR5mxrHEmRMFU8uiqDUcCnUZjd9uP2K353gD0nfqUY
UE6Ic1XOqDUoS04A7ulzXn0R9skyQ/GrNSXyvSGhxPayLCly08mJTmmFkrJDBwD6D1w5HdyH07u+
+NdVWiSseEOhtYifUz2mULnq2SHIygDyqOqvpAiAs+YyGkXGAHZbEbwjy49PFUL5vc5c5pcPLnuQ
n/0twGf1s2VIP7TKurxW7CzOCWrdy2S90887r1Sp31hP5zrjgCnXnsyTQUNSjZ+usCGnDygGCetg
iTt5EUUNWKvTk5YntTHG6Pqq5Jb75ulA+eRfQZJ5oozTgMl+ax+UTJdhu2WuIkXjQLVgbTXGwQ1H
C4tPvqB6j4ipQecDg0PJP7MgbzLBs16k1w9F/xlq4zgXIPX6eH/7R+/aKBY3gTuBHcHCgEgSOs2z
pN16mmf0VxqdbaE3TxtXIb5kkuFee5f8wnP3Pfglxu3iOa5f7+u7UGNFCJbPvXYHNZjIiJ2KmrE+
coRSdF6LkwQ3qWTTGIgmYMBmK/CUMuHHP/vC4qCI1A36pGEslYwtqrT4PtLks5MVws0267XPnV23
O0oNNJGfR3l/yajrT04BFggMLk/bah74VSlpBm6d/t9v60h/1WuP6zlm9oAhBh+HQd9juoZ01Bzt
j/bG1zrKEEPMuhxS910weqMaLEohUFVt/520EsnPjyN9nAseHDTtHv9eUgmUb/tqQ6X5jITVE9eY
+7W7YsNhyBfDz8oRwUFvqi++DO/coqY4G7V1wnRkfWAqcwNvngvGHOuviN4ntssAA1OWPL+kLAD3
d09WqGdDBTyRVBk7p974F+bbBgy1BPp/BzDQodwAqbEP/yK5ynAcDuYXtiaMsEksvDloyTpLrjpS
03KlatY0UaA23aPuVJdLeXxETp0+ALZ0Oj5GV2KdVddNBkVpkuEWW6XyVn9JkjUiP3HiNwGdtvu3
QdizY7ThTJQ3jHOIa6IQ0kGVtqsBwYCMrGk0onjjbxKFSsjp9N0oYKdwbRAyY91pmo4B/Spj/lkx
2rk8UFpnacx93GhfPHmsAfI9Qtk2JBal2EtI1CyIzS/QA9qLUVWqzx6zxCFj7pV2tlxXU/nF0JAV
G0+ZIOz59pa+PlYRKZpu4Z5dG3Rj3rx1kqpbxzEx+MgATVLXMdVoFgu0kGEq1ctocxjTnhgrjrSm
J7wJBiBMDB0hUDpfPQv8k1ugRAQBmZXD/dZVTzTd71LgB/XfSmWHzIt69jm6avbGuIfPrmW3KA0J
6iAYU3D1wiqUGuh4bPoBpEfrb5V2X2kw+jNY5uYHBCCuuH2D8hRndic66/Dinlxv0WtLjztvdzkC
c2y3OkEOyrBQzNLeV4rsg83pJ6XQL3gZ1TrzqRdwZsLVBU3pBg2w9bSMGEQcGw/c+mqJvdbFjJQw
NXOsapop+K/HNDlw/5bgBNxJsTWPdYNjhKrx61srYnZ5lzk5rKNmju419gqDLHRTtY8i2KB822iW
BkKl4xIA485rVEDZcN68QhpR63MmyPOj2MwxyspEAL6tLWNiZ+3Ho2NclMHppuBD8QNK+gxmsnXO
4PJidKquek1DlenWbuZO+Kqi9kUsDR6KI1Vy9uYYuuGaOuF2SqOZGdssk3Hbi8Pz0OE+7yre09cw
wVenNLvWh2Ahd4Ka2wOOqhRvVbP3wxNZlk7GRhGcZ/fIzrWV7IRt1hhYvySE4LbbMmDTW6R3u7Qw
w/+b/ES6WH5mQdhC/OZo3jn9wId/+8Em+eWzmWF4Pph2X1ebr5t/j2XmclCA5qaMgxsJFAMOdeP1
bHBhpzlxqHv6ZGC6o4IHTS93mHHAFOXSSewtcn4+SPaEr/o+1pXJZoMBlXRoN9K88BDlYC3/9Boa
QK1vujhLAnr1pJHwmQ5G7pr8BPeCU0p8d1jEaLBMa5FLwaGCUz8qMtMtBk6LdxQ4BOcLjjiyrvCv
a34bP8BtJNK/aYCa89/tkLyVB7fj/kL1zLqZ4/F5/+vWfEJ7Br/g4j9W1TSrHSpQiIvhVBqlHez/
Axnj4RCsG0ZZwxoyFJ5Wd4UzwqG/51Y4GLt5NJPn1bz0bAJNzgVtLeLwTEu0bhHQf4qg3Glwsomk
WLoUtaA+cD8pw+0chxLd1BuxBJ5aO4pAwuFjSdqihakpF14B6TP9MW+0ELw197n+N1xX+qOvmEui
eZkk8wP4TNsupeMz5dNVI0MS/rju7Yj5CyJ0AJRiN+gNeo1MShpY08KDc18Tzu8lIXzBNQg3zG/2
tql/t8JW3CLhaRZWhgXGVROOKtk2C7BxGCKeruvMsSdbG8MupLU1HY7p9ZboAKnS0RYevdFb6nXU
CBE+TQsOWHFOsUrgrIsywy/kiXZxEEWTSueM9Iao7sl1G8KQ/cXHVWQzsrcr+zxef/0PpCLS1PPe
aXlAOG20CaHGc5Zu0c2zYH35aoGAy6Wd/Ax3jQq7XWTnrYIm7SkCstKS3lPd34g5peXYg29ch5hX
6zk2riwUXMkPmtOPz5mSQ2gxZzdc1EPA725yKxa1OscTGdjP8AvzWP6P2Av8RY0OQluwO3DlRM/U
fea/BIGILSfrg71n28f6pZ4byzQyCfgc+0QedANvpcmp1eT/BD3o4W6rwCI3oEYtI0SSGzx8HTUv
VQEc5KiYICOaFqIghQRv0GGqfPP97Mvh/oYAU9SWqGi6Ad4Is7fdKGcg9Pg7GCiZc8WmjAygBW3E
Yhw8iD8JLFH/g8Gi01KaLK4WLeXcGSobf0GgkKbl+SpVOMTiN1fwH0NeAHyPKmkzKnASVna13u6a
1zrtydPX5xJaAq9cuEOVD3ek2gGX/SdWouJBW+I2seBXOU7pjb6GtJ5Ea1kNiEZOgxPbuSYmQjRp
xn9BQKRCPMU60fchaaUGrgx+jXlISFlQ/dUFYkYWXgx/ZiX9mOwZ9T96uhiNpl9B2QoeNO+hmmuJ
FAroEzdCzcwiXD2Jeyv7AsNh/YtY5w6JAjBnTMquVMUqMQWpNVCqQa/tB+DvSstHkT/qrJ7fPGYc
3lDH9nOnBCAceC3estRBotFE3yvMvxYS6knTJLX5YxkuKwiQVAFn0JjFOzJ4ieWREFKdHKibM5cC
rcP5ZvEbX57Q3v4BO+0ZPXmlOluQQ4LJqANGlFZzyntxd2Z1gCxlEerCgNAzB42G3w0bzpdVX9pH
WLVrGF1umFhh2ycGU/ydJMPqfuHoORvwXqKxTpnqqWSdc1onCoSw7o/LtaAt/0+wRYes8q29blzI
Xk4Jg4BWeCEPyhtdfn9c3rxboH80g59ag9YGRP/J/HdiPBDS8lp6SXr3hbxkYMe1ZB0ViMbWKeUo
rrMhKv3ygFqdlysl2lsSEaduVq8hrP4OnU2WXdBC4Ce2zpOA9NNLfINJ/i9PIMXl2IfvzGm64yae
PxaBMJNKgAZyw6OU1y0Sn3y6/EHCIW/ZPeUynU2TLdqGloxdhw3+cccLf3iIVPH4znnpye2Jk4hM
Ym6gWVSU3ZFRoinUFJCrMWeJBuCnbucg+FoyZPcZMEKjdSiTJLpmXV9fLGyKqeu09ajBM67aX4KJ
auVmXEsDR+54DIV4LTxcYe5IZY1nGAZKN6nlCJ/jnbsZot5Lb2+tTpPcJ/A2MpyHc7ff7KOspyy5
rNM9CallbMkE5lNqG0hNg+DX975CzsQKRg01U6JJSSvS+ImPYAUxnxg0SUvIl9icarSWa/Keu+jL
W84FjPxAca6/S9IXtlA32JLxYGu+RL56mIG5bUyTWnvwfqVhQz8LJWtabP7Ce0yCwlliXcBY3g1g
nmPmlpZ3NrMI6BrlQTCW77qU3xU8Fr5yP9yQ1AnPLGY2AWx4NmZbht+2ICYDtzKpz4/F7+fWGCLf
WSRznKEuYlZkqjTvIgYxrimrCLzMVxVeytYsMZqUpYU9DizPkqBXfMh3yfavjOxHxQarhtNXaRu7
yrizooLTsUMpy7v6qd+3aNeXp5wTkEZG5nKhtj6U6BKJlxjdgiy+Yh5siFnUKrtGyDVsX8jqxypt
wrRZlp23AanX1q7loNPRqh3Jdbhp9WjM0G+uAshnrGKEyNxGTIbc5J3g9iwBDKp0zXD/9g7CKCjn
4u+GUJOaACo4zDJGsM/AHcctXG94KySlVsP7esowaWp8LmTRHUU56inN8lSBEQI1gSOC8Ccigqio
tJ4ou/QSfxcEiESrR8XoZhVbLBi9wIdnqeK7Ng+A/VqK7i2nHgQYFPHt3hTfi5XX0D4PcYRPhF+j
qEqJWYI95NZFJ55ZWDfJ3GL0FSY02+xgmDlluiwVqfUhNET/18YxtarQyqjaSg+/T2a/Q9UJZH49
RpZ8AiwkucWO0z7fAkfKB4pOtFLAGhILx4woWFoWFuSi+/52t/hjyZfbMXyHTeEmw8B3CzCYTqhD
g4dO9+SKpJttdajwxosYuwUb1uw/gRYVxrw64hLn4M+cCI9aXObad3ne8M9NoChmBE47lZII/yNg
9BFG9jmNFdoERjHUWzQxwJetVVFKWJ1LpiqTxbHgpDpxJN6VgU1iUPPhzHvVj7FCZ1T7SovAkKYZ
eXuagQcT4ufskK5oSAYmpi7TEtzBHmJEDMBOszFKXMLBExRSlWqqrieK6XaCrtLJcHBhumn2KTwq
z+bfXp8uV2OaWClgDlwrfTPw0LlHCrYHuFYcC8kceCNQSfTeRwIoGdiz/sCDQKCnyf9JutfjF4qr
JaOGT5ZLIFqxwFYIUDPuc28DJNhmm5ryRKTrofxiV2mwGbN4kOKI74pY0jIJaFTBgrHjyuazfcjv
GvBV1nQeui4NUkXZCQqOB7uAQTjcjx7rhQGK+t4+GZTkJKA7ql5lQ7XMK44jQIg/DJ5D9X74zqTi
4hkf+61JJ0L188Mxeg6NzXULV+pKpA22xWW/Q3PKzrhRN9T6eUl+0N4XcrdBMKtgUHVK9IbKs+4s
DBD057uHOy141CcmblHIHrv/BqKK7+JVFPYxJlLJoSfsEJVfNIbhKPxSq3wsa5vmbl5foj0s9D4G
hEtEOQRktpqOAw4nJ+EcTchbljYYlQpqpcKIQIV+XIE0aQWyXRcp1Co+Jb+iSj8Q4xtOJwqz4NAK
NyU66/YfXdu+rQolcWTqoO5BGohajG5sapJ0Mpnvvtyo+nnKYlkz4weJQ5Hbjvxl5oDS7tfwVWnv
wsQk5e5lio5lwuWd7E/6oCwSnu6HSm7Qtf3hOQDAPPFES9GYxVRWWSot8nvJAcQHILG7iQlzo/yP
I7+J8SvG3n2Jjm0EQycabABiKFMNsPPXYZIQ31AlfplN4YxbGvGV/CaeHjlRgTF+OxqfzIAMxxz4
wm4+6LIgS3C1araFjhwENgXnpWEDEAT0kdO2hBPTyuKUO6sWztU0K0bCmO0ppAp0e/141ZgY4BdB
FFOWSd/APUg9+cpiu16FiYOuvQKPudI8RuarSH/j0wc+IGCDRFlTP87hBOhB7dGJPDgUk1qjT9w+
NTVvMaiduCD4snbG03/bZQjHwB6kd7GKHAgqf+H7IiivhAPYSQntU3HAHemy3mhdYTRcq8eMhFD2
YC6zAHJQkW2VsR3SQwzuTa2io3LKgfqf43MfTJYcpOWvjS4eZYk2hy1rffcIN4zl/eJkbIl34v6G
qKG9dYRvrcDNpBqa05qlDKGxkhScBcczBsOdYQ6d8UmiS85JJEMzqgzhrhanx0MgK2dAq1BhqkKm
iWm21uwiOx659529U86CATwfMzg1A9eF0uW5j0gvb/lihMjBHgu8MzQztva4lsxCqTFdR2fr5Utf
TU33I/89pUDXSEVZju6p43+bJR/edJg7mynH86NUeYZvXqLQyiOoL5h/H9/ds0zQF2DqM+AHE3St
7giZe21DHvL0yoo11k3XWVI3zZR39BYcdcQLOqEY9riOH7F2ofd4t8Id4Co+AOnKN8FaqHOvGYfm
hUfUYYZiaw/MgxOGNC4h8zcZP+zMEZw2j1OsnpJjaf3uaWAbq+UEEeSWQsjaJOhj82JhZ8ak21K7
/1651x1WWFrM9Yy/v2yLPKvt9cqg8Wy7tEF66dO8VtCTdT5LkqaGEkWYEBWhGKSaF+YEyVhsW8qu
aBYfiAPc7MScomIOcDFev5lP4NApluX24Oexi2qmUhuhBWSJey24hNaO2sg8ttSbf6lwwrAWi8Wa
27jilJ1vtLTYpN/k+o9jnKz/KuGWShrq/+ZjB36wXCVXJPNffzE1sgJdYaLs64jjI/rJZJkbnExP
Ay/v4IlyOsZO5TnQK1Sq+4OUau/XrJS5zdV2yTPG1H37r5NIUVjLn6wcODKHW3gxo2YfISauyY1e
ZxH3jpChh8q9UUMEUgUvEdhtuAt3bSvKKOQ4NFZJI2wPitzGkdtKjIkyI0p/b4n8wDaDOENg5cCD
eSmYzA1pOdvW1qfQcBaKkXdeBv13hlSXgCmJ1fhDnanukROTdsd/aYR+35RI0E8hvlreMXUAJ7Ai
5IrMLlad4RyuIMt2QNGlASOVfkuwwoRMFg78EFQgio12Jbx8bUuagcULPHarvrlaLvWXDR3oTUW+
8DiAkFNptwKQieLsxbqCCmuDMFJR63SDRu2Q38GDDg6yJF1w79mLPEG2nFlMiNJvo+9Txw+9bCYC
28te6y9X7S/64UZypdwEfJaHjX9VVRYZPyx570LesC2snWUNqwma4d3I3ahofMKZC1eTVnX28lOA
xM+GzykEnXYAYDDLhG9eYi4Ws+5QuV5iMk0dDDRkKehh4ILibZyydx5Q6CcuGo7yYANPrSNP62va
6T5s7tqRARwBMvjop9nFRzul8hbU7cSOljB29MqE1nj9TzNRIJ7ZNOuWYqmt14Jdeob0YjC/0BjP
bzQMzVP+VoAeuORtPeHRfYx8A+Dy+WE9HbKuiwg5yo8nX5qv6TZdThctwN0tRQcUpXx2GmouUu9F
a4Dwxb/hHXZlALfMkCb5N2wdT3w2J8NubGm2sAd4tkPXh3L8BagzuMiEesDMuYf1DtXr7z4IonUf
79drSpJ67egeDnhBxszfIYLO/kw/vYpXleQkic/aWHQJ12zw06TCYRig4kZho/WsDb7iEBnAJjI+
TKZDdDtKGJE8P6SK5KNJ0ua3viB/lnErG3Eo8CbILzRF+wQ4fPdhRBfJSqMZSXtlZkaPX3pPfBk1
wJYlm5rArlVX5iqzdX29Q8l0NVUfS29pn/FV4nViI68cv/nCjBHKR1TPjpVNOlmDFijFS8/9+Bb8
vHnThL4fRKv781dFrCBKQY1mG8xGHcrVawI2Cz6WyDA5o9Stm9AUfVEeGReAUlaJlyGIEY5xeITG
+/lQ8B+yp4csGHzSPVDLOTfXUiPZKB7zKH4PHdo/kpQjDYXYWZZeW/fyL2bw4Xv38eFqkiTz0tNR
vBO0qmI4dcmiSQfreUlt9lbye7TH+WgPYGeBc4co+3ibQB2lYsM1PNc4LPSLNTgW0QwAQxfUgK2n
rtwWQlEhW+Z8AGvUb1b8KeRKYNLYCiLvqpN5ky22aFgT964y0OnpFa6jaZf3RMu8gKzecDyqnJMH
yumNpi+uDEmAnh0v3JyUxwZGwFfD5o4KExG22wmgdNx0dvHEEWbtNYRwsX2vIvfVmyg7YHtmOZtG
QpIbqU0TnELfd1twPIadFNthe7BHklOsO6pEtnY4A87AzqXOZPlXq1bVTV8Ii+SAMz2Jfxt3SSWY
h4hqULymCzgnZPJ+avaq8jwUiX45fP2O/v/veVYKbC5cx/Qk699JfI8Bt32X5FElGiXOjxQtzavK
zSVrrB1UmSyW+0TTzpAxnK+gq+DWHf3uF87JOn70TeaexEgPC/nUkOxPappPREDFqcoeQTLbtMeA
AmHGdHhiRObm24S31vZEgCd95I9ZqDVUxJg9JflQ2AqRPs+QQYnczxyIJqngLQSbxrCJlBji3x9Y
8ptI7jxGqaBWGDwYKLY7+nfmc7fGobSKasvSSGUmGztdbkTARNfcpxxyQA03zNpVLSArzegRGEHm
w+nCMm5+uAG9B4lQVfgVpBQLMv8IK+pA1QE9zAbHk4AWTh6nhqF9DfBHpRiHFNMJSL/gdi63E/AG
Xqq+/xyhk0wVuG2DFG2KvTAbDKySJ4gLd1Vr2ODvogY/fzAESXXmi93rha+rYc9M4/xiMUlF3AKM
oNpknpCW/0YiUssJg6nOwnt9R0HljnouPTCwmtOe1EjIOBCn2Y0pkJWptmbZ2WgJReVtQHhAzAJb
fhkIfMD65/Mw/xafqFZy4zfnQNJuXIgQhXSIp08iRGceLCOohfuLDSKWmYWI5twXfG08E2mzGNMl
XYjiJYjouCDOmZcwsutAtkROx/BKL1sDK6nf1fWdoKYQ4VsYg9uFeveDpNLGraOTavskCZgAU1Mv
1pZC6AQN7ah6s5/8RJjfdpCoHTH5+qQIos82rV+d2Af8jBMO/Wl/3WnVtE0tf4UKql++8FbLZIRR
Vqb4TugsE0axsyGWeGBrnruy/IpmbCyhmQpcD++Uds305PFgCTTYOSJ8q1aYdPLMysKUKM95B87r
wlSZ0J20KZ61NHS19sH1I+ofs3V+/oB/uiF8TAUJ2TdU3XUhMtfx+ZKI6lXI1mRerBcR0GmW26fA
GMOFwkTYwEzOjTFzyq19b1fHYxCXegMIUcflx5uuUzCFD1k04l18Sv0fQQT+JszeQBpqwHjLr6L4
8GKmnUYAPjDd+3i960MGq9IEXj/1Cc1MxbB3UMjiTnGW7C7KEqN4pSzLo/ZD++Gc7Wn6Ffs/jTXZ
JgJ2IefHmR9FwlKDENNvkKZ1o9IhuqYmoyvMa9yzEjiOgbU38nHrjtoeEdJIIQSAESC99prb4HQi
op/eBsLrneFl5klLtu6cRIlvH9tf1AwyPN6prgHC3JOIJv56t/42sT3QjvfliRXC8silMUtNBaeI
eH9d5/s52rOiXAB6hlElXZvMGekB7AC+n1JgCKffLnIgpMShgoX+uWfpkpnUZgxn2plZxYlunG2s
Qzh/f3AC7Kp2mY95g4CyuSaGUp1VKvolAtUaVEOmWZbpbY8T4KGfji/kxg/jaAyeVESKX+jwHT/r
uFcYbGE41WBwCqsQ3gjeYRVxfUY9R4Ie8USLB14WleFGfB8Gi2H6265S6PaX+AjWWWPJthOSNvIt
WzHKq635UfW3GbevFJeZRMkt7uxdnyctj0lEZhD3bFeK9AARUZEjOE/Yk2Ikmry1wTcjC1DhqD+5
YNYDkW32uwxNSbw9i3mE8WKTcO5DxeYajFr4nInnfho9Q2zXDhMIQUwntE8dvnicUCyQWwkLdwZc
htLxTsRL8JLCsVkkOBcwrmWk+m+mw8tD0sta+AzeOW4uBwfNF9JXIMWRehC2g4nmS24lHsYbheuC
AR2vOSV837DgDA6JwjgmXb7PvtA0Rg0ibBJxdyPx5lGagoGAzz5moAE3OE23laWtpIADgFjo42oP
Vnkgxa6yofuX09vmwLDedgEmF6g8aDugE4ozBDgcfJsQ078W3I2WfSLZxeNbJQEajGuSza2vPSAO
H4A/F/wnC56m/0Jj1tNZaOhrFDwiFFQAQsud5Orv//h7/iuvmu73vKgMm+VEXesUYG/3c91/ytSz
0gUqGCTbUh46U+htZBgI7U3bhIkEbY7ERNLAy7f2bnS8N8x+FZ7nuV3wIJcfnzILNsdnNAbGEyrF
nYM239jtA4POsIEMUb4IfBbcEUc3uoWJeef7QFl5ET2N0tZY72w1gDmVZuWqlEgNc7W3DJMabbsH
tcEysdFzjd2wtCMo/Ja7nl7Ig9umepFNuvYE6G4ZQ6OFOwkyqeNsypD7Ftp+SHISYtSEVKG7VcbW
NzmCKdHTkKrlw/ZU2XOwUevTq85gWL5r7gacXmNZh3TLSehsF8NWHgL7lhcKOscCMqE7fwbFVciU
iU4KvsJ/yagkLEyjeeo08faEf2DjXDycTGmhLnKh+o9sA5Eys5cwAm+a8mHyTIYl2s+nILal3TiU
1qgsiPifJN5pcdDNKd0SDPEZJsnx7fAzhyGKCp375ElT6VM+kMNdMc2V0xkyaCEA1wDDOfwZ17Px
fCwcT21zq38UT8u8DccLPVRY7RbAWKIcRgu5NcGh/vi3QQbXceyUPVAUJmu2tKAATa/FHQCG1+k+
JZL80ZCe7rdEUNIilPlCjOP4PtztynMPDrBS1dtO0zLL8cG9nf7JtlsrNJI5yWc56h081uWS5Mif
elLmnstvwEjFebFOKiLv+72GyU+rFNkgXUjF/liR3D7n3P7EWJR5nYRkOXxaKsLQ0ytrB2hPiRJq
pyO2jyihQSEHWLSxhHhyxFdYY5ETNETRk6bORHxv9R8X7wNv8tJzGd7AiUmyhTwgk6P70T7Y0Zmz
7KqfsVb9rOtcXLzpxhltYByEMbcgMQhVNZPf3v+SbToKPvyKEV4oTDu7w54Bqurb3Txik7w42EII
I4X5FJkbSTnJ3SYioVXBG2IWdrZ70oWFidzp22ZOrpfe9zULDJ3d5FrGFEvNUIOoirNLASuNqxeW
7CFx4Nlx9VwHmcImW3MonAqw0CMAGhMWYq2/66ZoMrSfMiIItBuK5qkLnsKIFVV1SAO+0pkmxRDs
olj93jMYa7zt+99sCksE6CigDniYgskDrIYRD9l3jx3ZuOFHRVWZObcyJ5qGItVEjQuZsyRzcexf
+yF6QYcqnMFSd4JAjONaez4EfVpmfmZ4Xbbxwsk99P99WMTn5e2MXA6hMAfr0rF4dTrsUd0OImLp
PuvDmnKbPG+AwjlAx6Uvju3uU9hwkKSkcImwxWNs6yoEwUZSl9aR1bQ1DbbSbNFqKWeYSF5l62Sg
T9IlEdx+yYaY072gqwkqO49TwSVeEBntK3onNHRG8029KvW+SPztKzXD4TsrRjAli4cOL85k6qmM
R7HE0A3d3V+K7cDpO0Ifh4UUeuDk+04MbPU40cYIT+TuvMRapomLM4bQ8pXZyrowx02bWKB4fY7g
7RUly2c7Tr4j+gNC3uIIj2BNv8do9I0RjmGcrFF+Djq5evrvV75M6DOmIrOPdzF5vK2doVtWOQym
yF2CvzS28ss3cc1Camzm22B73DK5la1wMiRGw1u897FwwmqmOcxIt/0ZGvScHLuPitw/Mt7qZ51b
k/4fheOJDYnmLktl6tn16MyYIts6DhnszbRACaurtdvuWKiltSSpzj6O5+Gj2v1OH36wwU9anQjF
pqkSLB3bIIjFIx3C6d8YCLJZTjA/Wc8xz+0Obdg4ADP1r/VLeRqGXE1gQqQjPLPfsDz93BoBCOMV
7QyWCIotjfUgliVkTrfx2fNRC/B2WJEtF6kMKC7Z/R2vU852rHsP8ch/DXU+BtN/u8x7ahelqobN
1dXUYz5Jt7ZtqKrTJUgH+EadlzSe2Q9mxyFACZckeloRyILioV000b69zDssYOpCzvt2r78rMOKc
h7rf31gTnNiqmyA2X3Dct/qs/e5WhMe36tSRMmaJZqJgkhjJ1rGSOAPygsHJoofD/eVjwEp0m+J5
7ZfC5zrU4iK++vqO9YBIVkM3uXEes8ol2ZbbpEoSEkdcCS+ysB3nHjvbJmqzvhfeY2T/D2Q+cChY
VEmlskofhapfJ0GuCFDmKsfMqJYR6IeB462/CNj+ZWDKzIuj6uv0tvT/a3Cjz7qTMJK885QvFzY5
1dzFNoIaKWhKJ9oByUJlrw4Xm+BW2ppCQNprEZl8dzQ27irSKytsD6vPjBhOsApNAqnhv29rmh+o
4QFAMOTjmd7s3tJ6qWuRH5zWgHWDOaIlqQWxvxkJNTtg9RF87UZWeIyXtk27joz864fHyG62wRX2
epiDx4hT+m1Vru3LklBebayB6QqpgIPZDkyiyhbbKDuZgfuWGq8FFi3cnKdd91F5jIxiUVjQqe/0
Rv0n8aExjVbZxJ1QDF/D1lmPFIEtZ4GmtIbvRdaCMb8sv5Blh35l44m4F9MviqV1jUsfFaIdipb9
zmwaKSAjKsegvEIGp0Oif8unfOsryZMpunPOrLVdavRA6SgZtCppDB0UgEaxty/aEtQitjUc+Ctw
ipMX2/pLYDBd8/gaXubW3ynqV00Mkb64IDdnfI5nx0mG5eIMqAkSqwGARBEAviHto49LLd4eviiw
t9C+Ap7EsJ942REwJHMusfp6J70fXiV6KWmxXiwX1cUWRkt11KAUfj3HMwlobOe+24CS4zBHgMMa
HoA85bbWCG9Cx/aqk+osZLec98j55yaTIqd2aAcMOq0lCkMjkEY3N8d8GncHloliJvfDP9/0IJ8H
JDIh+blQ+zgfAAnsxIiy+Rdv/v94GrCihcbyU16HIQam0GV5tcPupCwsDH0fjhQy+rEImyD7VI4C
IIQ9ZldC+BGPT9yeQ5HxnvVSqCcIGBbsi01fYAPq8GLYb+O4bOIofssdWZjn4o2kRVILXOMxkyGV
AmjzG4Ojx+HFn/h5bQWPtejmeWzpJj8afIByv+jPiBtxDD/T0vboVk4B8oqVZclF5rTT7VyXYUz0
vo9qQhilfefBKfR7Lt4wZPk7HyrI63iNNiJ31HGLgeOedJBSbVK8+DmI8IV119PW3VijIMq/J9Xd
fotOTqFdhRBMfvJVz2RSaMU9UTmCtBlyuyeDkKzBxyD1AVb3myZsoBQ90Av9WBja5FYWrhGXkUY2
v+IDEYPuOKQsJYRvmW6IQdMeNgwYNYJNhaAxvCIbjltkqqFfmqerceyzpm6LCFyLEM9JzVKHCJlM
8zV5TLdPNPua2dYFjCACwIoaJthiJ4Meuh4qBSTdCcwPmUwYEz1N8nmyTu0NNspzi0jMwGNOI2rc
F94LwkFstboca2zBHzGvZ3oyzjIszUvxJTzizBnWYK7r80Cg2U4AHQFl/WOF8kpPY6ST+l/PWH4V
q6w7+A9ZqJX+EAh7coYIOHkMM3IPyWdWrgH6Mva0p547LfeeURkjfEfcCDQ9ZaICa02kiTa/XlNE
GN6AWUl+tgpVxy4qIUKtDI10cr0SpboIxrtIiGSPhS5F/ShzqBYqz37PapApS+tKEK0LqHbXRIG9
r1omIdqiNz0WGZes8d2dPWpFtwUYQ+/5FHQcD1SJzrPPj3yItrrSDc9rPpYcvD2m8yvpJQQldYtc
lBFFlyCeNoT7QVcYhcP2Dzz+0gxMCB+fbc5hdSaA99sKLQDUzoWzq5lzIDAsARnBUAKuUOwSOhNC
touFwDzMgwPh/+YuiZZqEgeE0G9z2QzhbSWlh/CN4LaHalLZPzLrRwBiBgOiD82N/y/6+eBr9og/
BGafH8NEA3vcHt2IqOB1ZiTtsOl8dIPK+Geml8I7El39BDq/vi/kj9OfUP1hKtqPWEDacmpwqlRJ
+MqPXHxMttB8UuH917BNKRoWzfmQQr0OsWtakSiTgDDic/bi8oSvEYpRvks2hnFabTSkuNA98nes
o4NYcWiXRjlgeXMJWQIAUna5GeogURtkwVwho6gQgZneWzH+ewKEGNORm5foKLzdf9a8LmcfDh3P
Kl5jozPrdREJRr088ohMcyK150xABk5vKdEctKmiJfdTO6Adx6c/98ceZhfnOHw+4gMcdGuTOdai
ki4+NBNwif6DPZ++4cCYqCXdyVCHKwICQYRff5s6wh0+qgTPDKyvUeuQobsj9q7MEuM7qn8TlG2W
Sy+uiWLhUGR3JcHgmhiQzw9dFuJ9oefi+cwTqm8smVAqGZ54AB48rECnLwZaSG1lUFCpdE+36Vnw
KJ+BnLb+FSLiFQdfgLIEPtDUai9sKdAv24Fbo0Pye0aQeiUtteUQ4sypJiPMfOGrJfhVyTQzOjS3
BZbwaallUTVbS+7strwgE4ImxPmfXypMyldtG7H+7nyWnmZgRkpXFxMpdRR7/kpzX7FUl7ZzO01S
6oSnPBXXVmnn7F/+Bz5OoZDUftdpRPs0gEWV54KwpZWieZ8RGcRPEj9kzNk86JyKqw9s5tLtHE+7
gbpxzbvx5hZdKCjucKA/VL6BQI2No991Hkj1MTY+DKkIu5b+CkMpPvHQ/vI00C0LpOV1dekwUkrZ
yjOyZ14mLgirOocLpttU2/Aiw3DrCSL4cvWrWiz5S0nrrxY2I4NdfATxS45OHR4Sefm7pyzzjJ7i
yTDPvCLjuo0SPoONxSPmajCfdf6ZdZcWhbm45xpr5tJYOTHl9y0gviZcIhq6bMpEvbiBfJ25EYhG
wwe8NB5ZQAihmaFWzWu3FjC0cMICfpebNR43ncl7QXSI+3a5x3vuJ1L6q0iNAdWgB0d5NelfLOoQ
ywwoqat0GZxPfwPbdOEXLq2qUrHR7hadp/Szez6KKOeCdf8Iot32rYlKwiZuZDKsfgLXUcZ7wVpc
A4gLdLaRehiOxbePzTN8Q3wcDDTAHg9CmegUy/2B0sNt7jXELayMenh8kaJn7uUlorJQ9KrrJsOw
UFwHb1MoScOWy4YIZPxz/fDOOT6AzwSn1MG9/5dC/6IACkBbMaAhyUAJh3+4aRVAVASB+PYhVyFx
T0iuzJslgAC/mX/AOwjW8sHHQDSIAMpF3BxLomhQBcCXkG+ZGT+fV5Ulcq5YxRqfnY8S06zcStQW
fmQP7uOkIlSatXF5oSqiNZAOWQYI4rUVzTDgXgN3RwDmrQj7HkBtYigW1cHJG/NSPk0y5gzG/ItE
o0mR6atZcQX0IGhg9QNChATuPZU6/rMPdAa5CAG1tVhLug4Upq/yb/vis9bmyKmDMW1+BNm2l/Yd
JCLKUgirJ1zZHq9FE2Anj0njf4FTjONK+nIGoKnzZWajbtxS3WmXoUIHAqixn+FbATDeqiHW9Xso
b+82jMGsTAovm6Q+CdWEreCIEId0rSSpou5bRzvx9CNQpOyTP/qouwDQ9a6BPM5OWpVwluvAaXU1
Ro+6c9S60etdq18kNsy41xn/1jEw0iBb2xGk3hJInU7W4bProotlc2crD3KhZy+WnoEw+Qkjkrpo
LRAJM2EwuBwve0gfbNfutD4fI3uHxCtYjur/5oLd6FoVvc5ePt7YsHnw8Km/dlT+78vjwUiceRIj
fIjoUQqHok5Ho5qZsbU0vOtVt/joR6i96bvwNJJKXujNZdOUlgdHd6IjNGW9NuY5ps8TjzUeVF1J
5Ftwy608VQTwD1VXuSlhHIH80aBPBrKP4ZdvWclyv63w1u/1s0GaB/YZy9r1h9MJgSs4bFo0V2Wb
d9/JmjKyKuUtVBt5yiYfD9i8HnbO0oMhSn/tu0BYh3vPVVkF1jQG5hjq5+qIcHjTVR8vgNq7rIa6
eRqO67NI4CDryU6VjnzVakjj0SmQ4KGUqtBryT9zcIb1Puc8ZNztOABYC+6uIbI7hkogsgVkwWw5
IIeyrlS1mAvOgUW9QhF2rkP7IPyEtANM3SKEUnd+nUWp0+S1IYCnSPKueqQ59jakz0SCWboDhtEr
Q7MutIXbMIajq1eZFC3FA+KrAOKrk7p3DhVYrxVWsMFKZoCAxe2KYFRdYMx765SPk5zyeGTTsQY2
7zK05JLUkeK0RkeVOxyrzxPz6OTZXeRGmhE+z1OrmGOijDXHE5jnOidYKV7DQ5ej4SEOVashPvO7
saW1HDg8ZFz2B9y4g7i97Z8WRxMWAjF+2jivUkl0ZfZC2SZxJ2LVAjZKbHoU6IPHxj548DHg+p5T
as2tOxmrLVgoDlGL1dgcFeRUPz5+PfozF+1auMmy8ER9P/5Miw5fSLn415BWc4+ql5ER01A2wNAN
abeYllVN5uOxeTpZEfj+0SrtembNjTrGzZ9msSNeQ0DMGN7+j6X2v5NpNzm7vPGGhR6GYeVH+s3D
mEBXzVweq4P9scLzVPHezDh04ykZeSvAhR/4CXpmPZ+ONo6qgcUpnBEAyG2ghtgwFtFodjpiacm9
t0jiErsf8g1B85urZaWquhCtmNtPP2uK3rOXL6anZY526vC6eeF5aCI8ElL+CwtrXp/kGEFnrQ+o
7WPJeQRTw8jC4AjYuO7O5pUBj5NLsjYr7iF5zOhoK1NgffMRi/sSG0LHy1P6IzpvNbkv/eaTdAYe
lZCFCtimllWz7XZfLl7mC5mEmX4ZBnLvj/ndW9nj0yQ3FVvcsF24D8UgGMZ/BscXlot+6oT3PNBA
rYbco6ZiW6XOKPNp3/KXSsOozrnqnTCkYM+iuamPLL0NEiylnoTTvtzszvUCpvSKY4bnvcR0OYiQ
IY5ENfpgcfSh4wQ5MIkR+uh7D1nDCJFjYJBVdrE79N/qoWp/GOupBmcMLjQi/sIY1KNte0lvhQ3u
Ta9zEu7KZ2fX7K1jIYB/8CTxeru5kcSeGOgjxy27iclBusk/pJJqgAHc3YXzCXT3h8eSqFC9MqJE
1brAe/RqkBNOrmPvgcuJwldaB/49/B7LaySqvzEaL/aduJn9EWyMrhYzFl5ZKMIl/tAE8/F0n0cw
agD2/cPQDTA4j0Ts/DGaqsQbmxknpZ49ccdHMaxw+bH27cnKro00LDYcbjLOloipbmSF/IMKj/Nm
EoEqu0/wrI3+judwwVCdQiORVq3nIkGGZRmRDFd0hIE+pZsATdI3REQ8ND9SMzyZeQQ+n8uNG8v0
ggZ0ghxD/m+KSeRD0c3lBTH4AceV9JMKt1TJWP5RVtPnkiU0TFfhEwf06jb+F6UfCRQzwMW2+DSn
tFxQWG1lCP9bfVuzskLigMk7Z+V9tPHC0sIPmSZ/q0o13luMV1QAg9ibMJU32G2N6iytfGv78upy
o1meVsl60GQEfmBkcZkKPOjCv3FSrAqlMZ8yNkewzcAx+dy6kcJVKlapEinOQLi4Wx7ue+E0yz/e
ADtgq8ekocijUB+hDxBlNGLJJ5F3abnT2fR/d9agxlXdp8Uhc/1H3kU4n4mD5Bax75hQDROQiayX
hgK8HBK6Vv5oJCVsPXl/edInsx+J4HrIIhiW06vvnhyk+xDBkOSs+bzW2de0+3V+neY3/cwjj9Od
6XdoAW60kyuJu5ucYfyfNBqPeMDBuJfPna8Qcp7gtnWeNIRD70ZhxyrVHP8befHv4B+llqWiqmov
NYNnvuxDGE+JxDZrJJXWNbkwrri+pI3ZxiG9gi9ju6WP/ogQBcW3CdPxGih3AckG6iccImXaDrJN
py4A1bOWcUIW1VLjydzfJfqpdR+/0Bmn6eaeUhGShQ3eyZ02hrGyW1hcagzEouRMK7Sq59EPFEXh
Qx1xN9JV+a3iEhtTfk6R/fktMuyEMc8B+eCO4NepF5vqh6nLlepolfP8vQaHPaIdMhhQmQucZxK6
WlCA45GQQgdrLOJbEGNQ1dqAqDWXtZ3EGk6bTV79KvDMn7DrU9tzxf//ilvhLGRUOzl4onMeZAqn
A0UkExO/PgaiS6PzbNSTTXBeUsMC88VKgwj36faA3qIeku6W0iJ1ZxmXKXzuJBLnrQA0w0maq+FI
RmtPA3B91efJyjMdR5uEEIXiNlX/yLXLR9/gqp4OK4nv3rKKT7gTyrs5uHZKpzurb2BGXjAm9Dma
5/duBfATldWHoEbCrlVPsWesDEY2ar7bU5B63nqFvTw6WB77YSa7Wm+DatCjrFE4/jynCCbhX/6w
PQYWZBj+oZSUqMeDoci672mMu7EtEUl0mdj2q0F5zGh0VdAdwvILZhblpvgx1liQtmFbH556dWOD
iIvN+7+l4dfDNcCGNFnxuPIc1TVjFGPd8F4icSxL0bDeJXsKvv3gkgLgVpdWB9/YKLI6oPhgSSDf
rUqy6TMsqCezAmhFnRYS4jNyKaGuySGwVw9RsepCE+Gwgml0Z0Y/7tCyPoAtUG6JhD60f+cmhs2u
J9HnwUqc3rAZPbaSxwXoykcr7S6pBhbGih9H0R3JXucpAxyExE9JWSPLg+PeOJqPBD3zwAm48Fzu
1y01OKLbl1ct5lSSkYolWznFtenKxSvgu+5ZLqISQEO9qnz/tNbYdrqk0m8TU3Gd+kTeV+pH9Qsz
W3Wi0XhA4+MJXOWN/Xz/0Wh97VljlQmPNF8kseNXjUsrVAiunmukUJJwje18sOmubkNunYqAEv06
1VMP2e29syeaWmpoeyYvMi6ir/usDn53+0eedyyEsbR05P4W3hcDfbLZc8tsiOMA4cDP/4mdRZd8
SkpCMxe/7UjOSpVG9JfMYYa7h9lg3NHrVXU3VjgfcwyVF/kGFxpUIjE6zMlI5YZG/ATXoJ/pnBym
/cbN/1MeNK6e46Ljtxz1SSPU3h8MS8sK+Fx9ghiv619kB84QAwDbVgNCDDTHawWYliFVPuo/Q73f
1vJbgNLLZuS/aMSDQTWcghVTFkMtKtou7n7vAs59kYZKpCNDxNQR7NGv9wTQXUhMCF6rvrQ0ScQO
eNUkkYIEGoq8QcTEhAw42cxNzPpmPxDgrxJj50xxz4+OkaJiWvdCUrvH4497GTpRMtr8mkXnSnC4
YHy+V8SMf9KN8EyHp3PPuyrk+4u1x+EnZ0fWgUdFZBX7HNtNpKwbTil6ZmjFmluumrVs5SDoXEqZ
XzIchTH6lm1nrWJefBL77FrgpQsM30mjXZu/dW08aXQdq0xBjuzMqB3AfW4vBEXYz2te8PkJ+Sh7
/rUpUD3jLqHPesowLmfosTkFRbPxN27CC+N3slWdIrkOGVw8CxBZtmohJyeWCkBp6cmoeMXnKsaS
B0KytCRtM5iULwriGIJb4Joke9uYp/Eq19obZjHfLZmK7+DlDUANdjCL52oHVe/sB8sR4Ev86FZu
A1/1gWt5pTs9XZ7qKxB5vzAWz/hd0YT4m5Xv8BA2SW4ElE3DA932h6ckDrev+wXNvVTwotVIDKES
WkzLnmQS7RSszCW8uZWP5vO7+Z32yj4RSRtN+zWakRkLSzbirAIqlTunAq7dFTB5KbK1rufkPSPl
xOhh3rHVyMmoZPGImsMcmfjFk/3Yk+oTe83JQzOkYThw53uzPXNHsHoBzpxplukGNzJVPJR8CfEL
OJfcDE69f92LnbMCbKsjFqLNz5DHaaM+dtKLmEhCybh+IW0BGomSNEx0r0aip/2Gx/8A/wNMfMjD
25AaK68ApurHAZd6ydn3tSAgaCRPXlGZ+X5SUbh0fRain6vVLW8+pyAq0vWOBwSshZqR1PAR8uwR
LFV/Y0V/M1z7llaUEd3SJZvCjS2hqBWRfRZIKpVUO4Gylhz5hepy+LwVPSuCsb7FdcBp7sFfc7Vy
sI7f8uvIx/oid45XgMwhgB1FAvdTmm4i0uNHEHAtfEGgOKyRmlaIplK6SWkULgXgbuAN+kHHOxv1
1eLSR3W5Lq0aSHLvG9WN6xZgU8eTTtTTkZgMPMgjC1kvcc6pRtR/aRW44bHQocAIGVfjWaQt85q9
v/GMOG+s4zhCp1+FO4BJbUpjf13xyhu7RebNg53Dvi5vM3Y1yg29zt5UZ5yJKz4+m9eS2YNL90ps
00xv54Wdery8fc88G5XeIEM6ugf97F/cqUxNLR6vF1BBUw+ACIFECcHETFOKrgNSD3z9NGEs8h3k
scWPji1NlcmvpXL/esCilWVaHIse+sZXqsJp3LsrtfAbW51c2n2z3wyWpaIUxz6IoF+pvK8ytdf/
lash7N8Lv+5Ye4MN4Bn0T87V1nor5QPRH1TmC0OjWn282bjyJruwKDqEcIPp9k713p+pKVVwvwx9
Ntw1hz5CuH4zinB03J8sYVDDBspKrGexCIBj5dXdJLW44O/h63Y3f2YajzGqQPDQibTvIgrKWsv3
HUKsf5hDyCE8pig/CZ3Kez0TPD6G1pfaCRZwnnCDYC5zOkORRbxuH2EPu3ds2hv3krnkx9SuayEs
Lu/mOx86MUsIIBZrEj8XhEnj14GStfUyGd6KfnviBVYRmgXC4od0HUA5eHoUaBVtaJX/cf4gHWHx
GvN9j7ejyFRhxyyOIngUI/rDKDB54VuF305QwG3Xt79yH9aYKaIExrxBbnlBT6cYys6Dx5ZJk6Wc
2t8VTjUqHoNoHdSWkd3MdT0x7AukdvsF6KsBBPOj+YTHUrjha+G9dLbevvk4FEOan/k1efM2BOUF
8P+W4jybquYa56/JQZORLmrUOozZ1jIw41CD2MQlyI1t6KhXkDdLFQC9la3Fhpb9PJuBSttyYsYi
7/CuUZWscSa6TFS96HbJNTjdAvdOsPdCGOKxofVWG6K3Yh6updmSH3ASSNTQvclP5bWYTrjAT2/H
s9Bi2b2kQAQeiHrPC90BAOybs8vNxPOQB+qMMcO5JxtqtqRs45ZhQspVq24c+FXljkSH3mZY330S
EawiU+H7vYN0wbC29mUs0Z+tx7PxSbiz1NSZVED2nwzOpiDBcB88Rn9a6+07sHCJL+0M+tnrfHma
JCQRjxtH5jsG2tp78SDGETsNLNWfmKlM+y6o7/WDP9Wi9yQeNm4XfU3jMVRDfM9Fi/9SEC+OqIGV
ytmD/XQRf9zD/830K1Uxb/CB+iWlpEyA/mUbNnjHCvtCWWGuV/8inS0PzSmRO7528NKf5t6QMuQm
kbFQxj4OQuKaA6P/l+5byRElX90CfdyWvTC1GeUyM4E8UXmfu1OJh9MeRtyXw3uYtc9ECy1Bs+6Y
2JYQ/ItlHjzq2NKiwLaLEkVc5UlFyV12E9wcjvlLnhyvm86gHm4wdJHwxNdpwmyxHOjN4RWoiSjS
hx2cBeX9uIEXsIJIrUIf/KFUphk1vA4KP60M5UNtDK9PVzLxIlsNGIGJ9z7LmegrCi0ZGQu7UBiD
HjjO5tms5OQdLk1HaH/HShnao7Z/FLWzl5Zf014cVHBe48SRHJpy6BOUruy+P2wmTLR7c5ZitSrh
HZPZfmBAny8sba6OnqO81tMWOzD+EHsGgwe2iK56ZGenNxsfvajhTJC9WvUbHn1MCEXUf7lLMM1J
dW759RoEiFt/tBM2aPMyIGk45iRyz4oLfv4vQRHMBlWimLEjrDH3wUv3R5UdN3mi2+9R0orQvDnW
KOChw1E8DrTcWLDjrS6KdeilZPe4fdTMKgqXej3Wo5B0FSwO9IVGwCoT29QU/51akmC1O1yICf01
X0o0cpZxAQmJdSWpxAO4h67ovLh9pBxmCTeIjx2L2OJNrirP7x8kX7xK2Drw5OwKOMvaSmG7w2YE
zBCaQuinEORLQdm3EApfwk22Li8pDdLhcYDwXrfXnuOpVtDjpa4Hiur8eIqiZMhpXBHMjBbr+aRT
Aq1qBgUY6XQSWLSKyijAoDlDsZBvxkuwSmpf8Gy5DX7AJDnS84L/yXe3VlMDeLHXE71TqjmIOh2S
fwiksmJnZRPDqHVJ0AdioLQYGCdGSJtPqEHX9XU9Dsgpgq2PGbtzMBSMQIJaU7HQ63SvsYDLm9yW
49uK2hcytfe7Icnn8rBDrf4fpUsYfX7kZoQp8mERrcQZhMMwkapE7EdRXoO0HDlexsZZNTQQCX8W
5v89HJHLkSAVXgbibVXyGGrEPh0T4Z/4H8D6xTUBNiDZNsSUQNNSd5Y4l73H2reHAf75OEJc5os1
83pATC4XOvIe/AQ8glthLTRQNcfQloFcvNwfd4dyy2Yf6WGRqi8NAVUYAEcpt4OBi3xGz2Plh+mU
Yx7A46oBC57g2CKwXfA4JYI739wtKQriANtROYuSXiVin17/pO9CL/tHrEg0SMpXatfW1v9H1JCg
/Gx+oWiPSt2cbywskMcCL/6rb+FvhR/zRuMfEZyuvfKfuWQpo/mSuYtfjnZYrnKGP2OBA2Qma9hS
yFth4zBbys/oCTrdDG0xRoGj5yFmGkZnk+FtIbH7zQgjVZ3KilMKrFkuE8iq69m36Ro8l0KRokQo
Wl7ChYLcAh3GKI/ChVC8Ju2CUhEW38FflV8n3Aqa/gOR1vDlurkhOhnf+vYlPWJ58EOBuZw1ocj/
hlfuOyXr165al+rlAm4XCxAgeWQinjgPhgM+NIzFLveun8StnvkjaQY8do3gC8whghxEbY7DHhH3
5NhGMgVvvi4iqp9wNKBLJjfx2f+MCMPZ5pnieXwTl/eBj3vmRMm0P6V3IeRyJzIbRB1srndRKy0v
nirkPz8f5m3hi7HRHA/AJ8xpQyTPvSS9rb2l2/4+ODkoRcp8qsH0eWXiQzvigA2hXcj9e31Horx4
sce2dUO0CfSspGTlQ9PLSEgb+lmZT6pSuV6mPlIEfnUBKwq0W0fZBIhlj2tJ5Hxw5mfIM/XcZx8i
femEPRvXiUVylrVcKkTbkpe2/Ikhgoz+YRc5Kym4Xw9m6MbeRH4Er0rONedye0g3XGVs4o7DQQbS
+Q/vSBI1bKddxtd52FOX5P565NhVDnH81B1hCyZyt0hbDlWTF+ny36SSDaw/8XiKLLlUtAw+X+OM
dARck/a+43FiXtODTZ3MbsbvSA8B5XGzUzKmCPMZLwg4vUQvCaotgjjCJ42qRESltkV+5wWO3EIX
2UgrQsXnUCwWgs3w3QcWDgKzgbmv/XnKG6vcYCf9pF2wYy6Q6QdhosQF2C+OsF9YTE19UF8c1Um9
nDrkq7b75wR3uDuj0yJMk864b+lSjhTTJdPPj3+FRATTd4z9r9w7vY7psnVJf5EBPDKEDrnyOMnh
hmZU9whoMLhgdQ3FEWcsJ/KpxFFZ76c0ppHLNK7viiRZJ8wP+Ln7byeAFx6hdTi4czIe3Ub1ysow
kMpTKv9LFvDfpqhCBrvvniPnuHa2/ICqZ2Kvm/y1HTvJjfd8hgxsuumLUvyJkrEfp5tgZN0whDHE
v/oP1igOGrew8wIGa3YWXSAIRk6Mfpy0SXHh7fD/oztFOpUijFJYyDi8NkbgvygggmArL6oDaV6Y
A4R1WKWkP/Y1QvQfoPGVmPQNPa6WHYW7611v/SXBnJfS14UMf271BTCvGDbmI4PTliNn2KSj4OG1
vLQwJXyFktXtJUdWrxg5mpZe3eNq3C5sHqzGdffYTDv/c27bqsb5BNHTfQOW/wvoAzN7XmwC3UkO
CmdVegeii0wzKG2DRnnkoycj5Y/WupgyOXIMGGP9zU7i2dD0kBb7hl2e+nFN7meDnjCbDnivqB+x
dZ3Q5iG4SQDKsQqet9iOSK0BkWXLnT3Rteenfk3SzhU2PNLLBnMDlGXUt1Hy4hCJQ2ook9hBJmvi
cohhldGKFpZjNXdldN0iWiC7/BuJGE+wn7zOiE6VgzadJz9l9mv1fbzIolcyIMxsw2I4gFIdkXW6
Qf5ewyNWkY6iM5PBdm6WPj8FiFOB8LZ0XpXAUD8A0xrG8/HhcypuMlv+pSOk3btQg+2zZViH+lMT
o3FYKPypDgMoFPHH/z2RthSofzcuJvu6DzWo4Z4WWTqvE1C9JXm9zhl6xhxRvv/mik5VKsiHoPO9
T8XjzAsFxAiDsBstE8QK27CmRbGYsNSY5KBA7kRv9E9LEfgYSXfbWlqTSqOwsUFiuuKwfKqSacfx
th9B/kwws7DKt1Fbk77Iqc3Nho11ehBUz/Kv6CtkI+OSuoUZgqbA8/3o3pdKLhsWgYD2iLgUm77A
1HBHF/HyM1I4KNtcXCOZhxdssOfmtYju8u7tlWnP/cdfLs7ZUbM4Av1kkud15PCrbhH9pov2jIbh
fZOaVYrbvElsbPAmA8d46ychqCzHUawM5qTU95gPc1A8moFn9nEouJG4vsWy4Z3FRv4sO5rs/T4H
VnDGSoFs6pXnyzW6o2igIzb9BlTEWRTr8FqugY8KcNyYEsJLs2GLB47EQUqwtrg2JpXnbI1IRs2D
kvjvl9WW7fg1+XQuY6Sykyh9Fw5AhxRV2+5RFQQDLwg77YjC0JK3A/rlIERYobcyolADx6/Pa1QD
v9R81zmKYv7fdaoPT109DQ4DroCl4AqFw36MGQouHm+IsrKGehzFJUxQxoiN2kSQ2VRxumUj4JZ8
9wNRb5owBeemDIQIS0q6k93AGzVhzZ6A5TzKr5R8OuRTnT07MbPJo4jnt+uF2dG7C5AuGkWPxDaF
G+52F/7ZE87SF/zGdX2+z4k7o9KEwNbQuEAJLEl4RKovOz2bTPsT8g1OCJLQxAnVDizCan1AqwBf
3zdfHVW8jD3N+XAc1cF820SFjasGGKdYVG+qVk4PLw4gU3sAHlsHAvkx9Lwtjo6XkljCoJqr8n4I
Yl2yr3/NT48uqeUw7QSsopBIrkwC2075J6aPFH4XWbLYbTpmvFtKp6aHwlRJMrjZ6OHEbEQGxMJQ
tR0nRNW5zDMBk0RdzzpkYn/d+leubhOjBx1oz1Tvpcj9a7RrNsFWxloMbTzDLkYjKafaP+dZ9sI3
T/xjyPW656kDPEooiu9ju9eMtiCZrrlYF1qgOvT5GgYe+A9WA0sR4VXqNaXpFPm5W/HKzXd4myoI
GEeXj18Med5n0f9Oi86E8enWo5kzPfGWo8+IF5z77VJamnJfm4CYWTZ4dEcd4sTXy4ib0MsaaGDn
QaOeiQikl5J/OVShxbYO6O7IttfP+wI21ZaTLF+UgVYrx2Zw3DpvzgYxTY67/YlHfRBZkt2mJARi
iMTJ0XuW6G0gF6vLl9b43L0Ye/5Yo+gLuxt7xvP4dZ9OA+/X71GWxAIzw4q/cnMr0m4Hvman4lPn
77m3IKC0qno3XSdJKW6UmEka9R2kWKzOyBrRewk0kkfOnG7hiSCCzNonanCm7ji4Cjye4DU5mLc7
dE/27io99/KfDT4aytAgwsS9GWWRfqDOGfOHZvskzbAu4UOUKrBoGIhmgKjSuS0aQYJekRx7woKR
ozxZvJ84GMi3J91aZ/D8JPUP7VWDa5LF0KdO5EdCfOoFvNJDIsBe/hAgQYxzvgWDqnPE7IWoU1pz
Toq94GBd6sKorRUz7Ab3uZnf3vxDVsX5bvO39dx8GFPDjbjtgJ53GOl3cOVIhw/g0v79Iz1BaIe0
8hD/7+UMKweziUeiVComt0XGpcHiijg4FDmsAJZXzT6ctApN9ZQGxzOWQATqbsV4N2aG+2W8MSUb
2Tkm6A2VGjMqRCmsgb0if78x58ZhC+riGo70D4/eR3OHPDD5DxIaUQjZl3xX3eHJjrFFhsfVuKea
QDnVBl2OUgPG21Ocs1hIbXkTTRWDmLjmmS6HHUC/YVbx1FoE50v7qJpyaAn3PH0xQcpga7ZwRR1H
tW78XtY2RcprMVzlS5bYz8beub6atbbnrfKf1WIvZ+HkW3Lp+6MvFBHjSZRi3lqtRh/7pcych5BL
iRksIZelHZkRfi7alLR72TTBgqZmf/9Xgc0/tf0xJUmnHpNqGhPhoVsYhTS+Vn96yjHqbyn28UiI
puaE6yGyRycDuSRO8EbO9EIg52AxFJ1pzeL0I5dQ37n/wjjHfKt5Jq7+YyGVPjfUvpiniXeg5nOi
ve7od0NBCQ3F5X+n1hZgdy92azWMGYF3O3yGUvQN7YgkfvsXflSKbxt3r6MQ17fy54Ep+fQKNRMW
FUTFgD1AbGnqfnxeYUnMQ1OvagajoAt95IrdteQgnpvjPM7dUrJoxLuyiSPK2uaRw8njjZXW62pC
p6x5Rd6nKXKOxkyEbvmE9/fLarVeMdhD/vHolk8SNnqLGT2I0RBfkwfpf/oSE7Oi/UGkV5AM4bGq
YPj14TSMalPkbEDAidabh7OKqqCEoIwrlJpN+0A9NEynEldGOaj6e8OBsP9B/mIIIVcv5I09G2aL
HorndKnWK3+nY0awV6t5IZMb5IH/iCp+gzBo5FC+Po3IfZrvwlhxGXrn0gh71mYvgPSBdROfCgSQ
bSZ/ZjwdMRrkqBya1YL1I335OVm2WuTroB3TeYh6taQT1kVIVLFwCtbzxiIvrrRWIZZOtoFYI7kX
aq4WwV+x0S0EZanHBuwEdBesZY+8VG6rvzL4Y694qI4X6C+wOeGu7q9st0FpHsQxNgLBXLWjuUpi
8JmI4Z+xYuNJYcDIMwnvxCZRh8x8ENbC0znfw3yrmDeJTbRZADzofLzxemPvLrCsq1k1+Hbp0jo+
NF9NdZyL/6853aWgEW5b0kKqLmzREQxOREeNzJ3jg6uuzHLHXKSa2S56OGVlFyCuwcJSHibAj7yR
zyHvj44ci3TNWJqRfvcVQanVo7ajCIqUWJyXf8OyXYzFD8tBOIL3mb1MuvwdzT6WdxaU34VIt1Fe
lPT3R/EfAu2Uj2aoyht5ttGSF5XQ8cCKX5A+d1o/RTGHlY2ALWqwRP1esU609I8p878iQ6alNWyD
tekxkxxLQVqp56Y4Chp/JzU06rL9MUZuqgh0a9bLYnGOpfbipU9R5WQ/HkJA2o3wxYTsn8v37hT4
TWgAfP9l9wtIovnD8xs3BgvVYi4hpm9VZC0d7GODDk8MksOYQk9DoNtdgLbuns+FA0Q9KmW5i18D
fvZLZpZLjxjQPtY0lAGsqXX7bf/aSiGeMlDWDBu1aW84QBGeV6/UNBObXQm7X7MdaU4agKdT4K3L
o/XOKUFzwQKAYPhaZVcqTJLhgyOP6XnxPU4Yj6zokud49D7f3fr5Y5JCA5AYqQYmD3K7OER8tks6
S/ktW/wV02iwoabuPkDGRpi0GfjvGy/czgT3J+t5dHxyEBndq0O5xSCCPNAnoZuBSGXzFap03XP3
/RRsqqcxZDB0ko3icCGfdhVWWJ1vHYa2MQ+5PagPRg3fHXbeGhTVvbyKepGF6qPGAw9um+AiiRSm
VC+BTR8paE+MyKlLv27+A6XykrAQM1mBZ6GpHj1nlPGVFHHgKm9I+cC+j0mbk9GvkVfVjyufeH0u
l83WsniYu5lP1rTdfysMYHt6hYb59x31AVyrF44VvsDxRNQq6FE9rabxoq7xbgzc3HSWqdUOdvuP
l+gnyF9rFOBKAeMp8TgOWBFD9GYJcK2VIHFp5CCeW2IdM00p2OvIk6QHrjojhYVFz5ho3Q/ylFmK
WymqnyJcF49OXvHwIX253nAIXSDJFFuWBSCSQj9JpNp61ebYYNWw43QAAHpmZutv/eUZeDXAZ7t0
2Ll8fG74yAfKajVIFfHquGgFmLnfmNPIRFwCmlXJWwXs49/BMhnO4dXEga8pgj9bWfn34QZCULEM
VY6PI0vBpepo2cg+9SaN3WVLQFKaq2ck8u2819GhSAPKPp6Uj9S1JRfgug/iNpTx8UfR/SRZ53cb
wQgYw1SBGc1fd7PqcNezQbrR5gtXCcLZtA4UXZXo+iUx6t+GMRZsB0eXanaLt7YnooiYDC/Ss16Z
r4DjoF9hwb2LFk8UKJn+OqoV23HxtVYSUoh3zlhTmAvcTVUYo9xCWdE51eNid5djJse7ClEExx1C
bh/6UShZ/aVCYSMccBTa7eofmtX+e7RIS0DZyvLAdsnFKBqV7ltO7WfkHwUW7APjYmNgkHivAlN2
AUe/y/BtiTsajAtYHLHQnVRxw1II5bU3//0LOs/6nu8J2DL5FBWZ1j59CNXbcSzi1h1F+sum63tP
5O8g8eCuebqCQmTQwY8JeUZczrdycAMLQPv6/m0bziHCy6SF8aMTa9tL3We4wuFZKxcAOzGkjcvf
4FSQRB4xegxkCsHtShMXci3PPiom0C6C9ZKmNIACODiez2GxRLiPL1x4Qe06hMtlc9kXi5Ievy45
sEw1Eac8VjhFrAsUA8Btr8kJ24FC/8IfQ72xY9gQfdiO9qSRB4GDhc4kaFUFJu+r32aMQ7OuonYH
6hWMCMP2M15PbLgMgQdyRC+UREx7h8u/Ipqfa/qsOOl1z/vLt9PmBHypjDnrcVrKGIA2GMaMXCFY
2TqtJ+efTHC8UpVgefYWl7Yym+asALh+7LDFjEINVXZg0+rJTumAWlSiNKB2CyFdwDOXhHHXnWNF
7GyPDnYyFCJDOCpEoFhbCon4GTX1GnzNKX8nA5DmJTTS8Qxr01ueEeAlFjjK0gSG+BaTIJOTiBBN
y3Bo/v1ufWG2oM4RS8hX/5VkyzLofmrimMWLBD0m8AihkcpcRu/qwrCxplkhP6LTSt/rOtil+PlH
PNf9rI0jBF6G1C1QwkEpFpMSMlDaO1MLCpxXnUv6BcdcmSlvTqwF2G+1IfOhz0zOqtLuDqlqiQ/1
AA6wh2iea/mfHzEkA/js9tdCEsE2voiL/cZbiaJalw4QpiAPiDaxvqNfa39yVsQibUuApFfe27BZ
VLpJIA07RZcmjxfFwggNepnXv0sB6yArpGFEGz4hT16a4Xiuu+egXyLnq+F65lhujRtLi8xkVs/v
NUNgUVBFDUSVqaGWoHbmfa6Il6955fxonFXbECVgskYPEHBuDWGsDMZFWtDvT1X1E8lTLv4gNHpv
5oNMugMckLonrs+JU2RfbqN5+i3ho1NyItl9LuSX4dWiKfHzBtioqiuC5LFgtwQWVCZRw8H8VvI9
yb92sHeoJdSeLrP2UMCPZWw2ObLjlOGNwM8zmtkVtxPbH827i8CiSuam0CEoakWwa+St9RwSwy4Z
XZ2Mc/4m7otiq9dRq3f9ndG+FcKXrDnGLDE+KEhiNcu7X669wfvidYfvwWBaCFSahWBORHMO2ReA
a2iEr7SmflOllVYxyOy4KJRM0anmfnF8GFevB+2+gtKbH1CppnnFLMgl6ONOFvkFHq7eUA1U4vaM
Q1W1P8kVSH42xUlC88MNn/Zpa9rfUdXvtHSQBREiJ9I+RqVZpYrkFUliAYJ7VcUaWwuEPko/R2nC
wrVQ3pvfBSy0TxoviZUNZIccohpFNdExNa77uLtJN9aulkrbMOrTs9rtGBPd8znCSz48BxqM4R/s
uo6u7QvZwN12+wSo28DUGePuYzkagWPcyDIjvBBt3nwhGsxufHlryErNbvmPpUGEplYADqfGZqjj
xTRl2wM3UnDu/AUnrTMxAcuPRUvAoOavzk8r+iieCbasfMcWail7xIdeVE3xLN+V5DSRxyvWZTUS
PlzC+BhxgO2xzRLP968N4sAgVM1B8KPxqoSvMdSz5Sc9gtj3ksd/bo3Hh/nsLPNoHLQSfhEQpWdT
VGufRpdi+SEG/gLFfqsw45mAe0RGDJ5jnUqO9Hw6C8OT/I7yReYqjVO9FEiXvUC0qJIh8Bo+OE4U
1YQ3xk2pvPbaoURGngSk5S2HkLpqsbT3WN5ZBc1zDdDM/oBf6Yqpg69qoQ4YN3/SGtvHoZdUcpQB
wFyDflqKlyvDNloAFIAwD+VOX9vmbrLV7PUPv3VMxz3zkC9DtqF4Lz9dsyK+e4j6dov3jf17NJP4
bU0zFD+m21kD1wZbG/WxoutdY+qR8jNXQ/OFZ9fOOevCoVV+BIwywA1vNzYEgT/zUKHKPXaTw1cl
SnKp0D9jS/ttEhbMRgYZyvPKxDaLcbyMXgD4p+I7ccw9E3RI4Clg8JiHIuikVunoJnMD9pUEyLXj
VUqgKUMTcbl4Ggh+wwcM/Vyok40/K3tOUx576dmtd7p3XQDSiypY3l2hrq6Pi6EhO2coVlyGjNpa
oWpcGetWESUGWjzcugo8tI3MATbEsW2Qpz+KGj8IoJS7N/NzxNqZZ6FCl5KNQ5yqIphBBAoVX/3A
eUg58vvTXTk6mmmxoqRZcTQHTltq1M5U7x5x5mzKDHreN++QmcL0FBoRvIVZ3gI5CYl5fCkmB3ci
1ZxBB8Clj963Aff8JHgIPLzyW756qLRD947HNeYExo8OCkWwNxZ5yesu6WCuF3TKf0HXgWWS5XDu
5LN/wUZXun4cBTOlCTWWbJgFsjVSf0UuZ2WGSZpYRdkEU22zCulbRDVJ9bU55e8qPLrlV3yD1KZ7
T/wNf04N7FGRTZ3SztZx1h/JkjnVc7EVMXa5qi4s5xj61ChT9rDxjBarn75zJFM9BQtNFD82hV9W
Ce3MMZWoXybkSffmmu2KEPU1tTI48ifKoUAFJYfML8eIFJ1BVqSJYBbpRid6oFRxW7/mwiI1V5Zu
Mh3StpQ+RDihsLJbwkl136hCNisLS5gkXFIZuyG/s3EmCEhwspspK/vsuJUeEKbbkGdCZETcJJQG
bxBmkAwc9pDnhqyDf6NZL0VpcDteOVKpCDiDpa/wLw1fIQaesvqlQS6xOkVmISq9tMiZjj78bGFn
DOVsCYD9D4vA4mDTqE24Sdl0Azu9iFfj1bi8X82q5nQ908wUMS0H2LfHD6vK/Q7n5HK74KxC3Kvq
2XTgSGBRN7VSsuzcm8YcSp62GyyEB+OHhBoiX+M4Y3j4LVUhF7Q5gtxswf1qaF9dY6N+9PQK1B9B
rLh7GdSuxFT9pDvGBd+tXRNE/o1OLo8Odn7tlxYit7xi9YrJ3cKxrJ8dXPEd6pwGFBLqDCieckI6
shfDeEL/0ptal4JE/0pni+RWpSHZ+OZ50WpP0vHzh3eRBxX/zzkEEjCvhH12g8q3iqAeQNnXE18L
jHHIjica3aaHPr21qIiLdioVmOvpEUuhPXTq2midGBBqF4Oxx+TeMTM9DcPcQosVf2yhw0zSUTs4
tJNUwj6GhuSNKsKjsw/gIrvuMA3pGOoMaYcgnxmvK6e8RiGj4plr7VFQRMAIUvzXHFqzpopcN9F/
LpjrQdG1LZEgfCm9i/4USKQuRORn0Lce4I8URWxmfFysiEB9AJDkhWlEsEcpTxtEllDC8oKSjeLo
Q/zgjog5hveo0DIsPdEt4irquWwlxwtFf2O9AMOSTQcKjo8FuTdbsv7HWc2oQdiSJ0eyUmkzJ2pc
mDgtw29Do9X/JiMLclTGt0cWDEXGSqDLBx4D5WXWqwlsYAS16WZ2ykQwqye7qDPQpNslUBXbw8KA
c5X3zp4oLEmzhsWS624NLEGGQQQAUFeg2xs/hu8pSySZLiLpJpUyNBvoUX3pCRa5iLRZ6Dlhc3ps
2A/8b9uTN+NCZyKHU5YyWW8X81g7+SmWDVfzmsfXsv9PkJcbMDFcXBBLcbqxfUSFideyl74IFvhd
cECqFE074PRz0HtmRZsA+7RAT5NgT61RXckL+r/2AtUA3mzv99kZMPrBpuQae3YhtpmH9TU6HrsP
NjzTNOZh8MMx7C67mAZRzbQvsGHMDIk/E/2wR2vIvBOdbCSFObBzpVLqx4u0HR+sAl632kl/PWTa
Y5pzrTGyAysXmd1wNYfw1ekFRaj64W1ioPf7wTUCQSAp7yHWUcTeOjQE8LsaAzPHyV2lwaYS5BNa
phpDjBxhF/zlUkXloNXJTWDRVvmOP8SCyiuaEvhypFGUsFWXPPxW7fVIHH5K5zdGg4INwpniS/GS
BLFa97cdykpoF7W3T28VwW/01CZmbcN+lfAFC8XtHpfbXXvIo7zWCM5BqzvvejIuaPbGVmUUfPVC
2C33Xvl1zGQBHImMLAxf6fUSTbWK0DgRovxaF3EP1MFG/fBEGqT1cCX3qbuhwdRis26oKuQ6FK8K
Tdm31NU5WT4TzaiKPjIXUz2meoWVi8Xc4+sO5eVnZ8/YVuMu7EREtHv0t4oFQ4KHrAIACVEtsYgk
kjrew0cTE/05f/cDUDUGnXVGgwQzdW4hnoSc07UmkcSZv511pxkeAw322tT+eOuhZG7mgy4dTKQn
cyrBAH7uQojboObHkoVgHi8IyiwbejGth2Z3PazCee8gMkzYLMVT0lVSwQsf6F7yoUVrOu+5yCca
Jhm6dV5Y+M2H48xLNa2+B8N+AYKL5zT186XZ74ib2wZkC5IHseaoI8AAfO1REpK90fNYOoZyLXz/
h+/SLs/lxipjAA79HBWqsSNtvjgNsdDe8W9/G0V5xtSis9PooGc0XGTFjCAHnalkBeAc8Y1DCXng
KBJt6ZHCwgqiKHg/EINi74/6UOoZmsrsAZM9/MZRNb6DpSuLK2iqQTi3OMIf3g7t5PC+hysSTNKv
h2rtw8Dc0MwawbT+Y5C9h38de4YBspCrw2QIkwxqkUaXVCaBQXWZ+1ubyW/IAvodf7Bz6kDcqoWz
REV6o8x7QKoA60LJhQE13mBPZT+3HoIRWjMfl2OPg7HD+0DKOEcjfzxWYM37IIAkQess1Pn14Ndd
+aSXsNHc6/Kgg9q/x5o/cjdOMLa1hILMvZLjRZ7BTlb6EqP+CZBLpBR7oSKoym5ge8OaRTarUHuz
+74x1/S0Uo2PKNRGO0VpMJmqrk4SZP2TI+LHsudWCodDvAyZjZsCJAVCv3WjUsllO3iR1hxOymd9
Z2FlqOkMIrp9lOdGomMTsQ8mBYpHJ65Kbvkbp78aBAMf43gfWjUZo5knmL0oqRFOwQ2pb8MDkrd/
z8P2cIu/17QHn5xy1Vb8RmIzDZhoqJPwHPahdfdeGalFqD6hiWgsAGyc/DLQR/SllX/DWESI/quz
80M4xHctw7OH9WR7gZK69/pyfaUz3rJsmNpDoW5brWpSg1/a+Qq9Z5kijPHs+lD+ReMvX+Fv6utg
NQcXFFeZqhRqlcRyO20FmCL2Blj/Z3QP9JlDRkZpHl9cwbot7jJm3jLlypzvcaWTnhTEMlg654Wb
T8p75YUOXZleo2n/YyUZnqQl3s9AwB3g3rDxIzyfBr086coJ2/bK7HKHgkOvJ7e1JvmBGYz4rorP
vrhZp6ah64fWgzOxET8KfucMxHug4Tgh4/YPDiShg9gfTW0vWP60gXpOsaySuN0/vNejNWnByjF3
B1lS62TuFGnwrQyDkd8YWy626rrOIfH2NcAfjuAWotfe0p9oHJEn/chEkIBiBwME4f5aJBzHFKmC
Dj1GHdjmoy4HfyYC4nnY/4tNAqOH3797bRHCKmOU8Mn3nTsX1LfpkbCf8DLEO9llGCIiVLEIMLX6
rryAl2PN5JhOR282o2ywngpSQdv/0D3i/fbAFGnEW5NSbdUNvGfrASuGIL4FdoiJoPzwKa5kRCDF
NqN9vFPdVVhO7jbt6N7tjw9DnXt2j5zNVu08vHzcuLMQu9yz2918iAFTnd82Ay0SPpFafGx94khG
po5TlCI9k1eknhQW9QqYUmC4iDfQYXAzJYKbjpBBUtKh3Wto6aYwjquDHeTPgZ2/kjkZkAbTZGG5
OxAYy1Dggry+heXlJARtq+i+3ikb/UfcvCigdILepDTmAIdgnDu6dEP/WWjSYopRe+EZ4zpLm/ex
bw9qqUE4hORZyku7Gdxb9+u34q25Co3Fi4XY3V3CfzeVi6BFb+Wf4XAHojudkiE7RB7QddhnhHpS
gTgcU+/GbxSAaHc8e1zXiGWLfekjwU7QNTJj+UIcFRRhwvKaZtdazlaK8ACpQLOUynJXVqeA7z4y
d9jd5cQX6H6YXEbiPzFgnTXA51IssqvU36Is/SjG58wS/8RlELwiBX/AcHSw+njqSmrB2YgPnxp+
+QR8RDygv8GkG8RgVWQTzMVFIkunHx4qOKHYAXzIhFHEyV+/B+cXm19caIw+ohXUxzZI8fUjsIRm
MvOrnFKMrR9wQ1tbd9IDBAwC20jpX5fyZN04pvsKDHyBPN0K7EWZAd/wIGSIXm5Wn5r92BqigMwB
OrjNVdk84YXLs47I5C8UvJDxwNZ5obkKWMuJ+NFZ6CYlHIQawLYGXOnFOed4lmsUa9iFNkxFFjpM
5MdOhqPJ8DCjkmbuIuYQYxiek/UjWjk184Z1HQdPF6KMLR2egNckM+IiOtYdsO1YFfgeyeP95G4o
Abxz/zr4wEw8r/AfrD9FBxX9TpgWC4h/7AVuUQCVEj7GyL87tZxQBvJCxYKCtD/4P//Tl011e94H
yAH0aEIqB8rSphAd18yUQK+7dOyoyYkFbkJUY2xbS58YYXEt7+6YCVt2L7+/fR0b2oRerh8nHypb
ZF+mneqtvH5iCYUPFXkbhYQGZbLc+vAhvcMgRclnR784VTbs2Cw8gD4bNeDN8tGCIYUlKSLbCDGD
RYIFk5reHX8u2gEI3kSh/A0okKJXU5uZxNrhH3hJ6/a4BsHeb/qwiRI/OZZvBFxteJmW7Fi9UbzU
ArnW8Z7fPVyea3qVXXTwuOo8QD6MWwkvKZrEyis1eGAAyUYLlWq9MdB2nUzLCSdM/bMRJ3jtII9p
HnhIvcCddxegnov/619yg5P7AvZkkONyGFNVmF9v/a6DyWi+uyNijWRjgJxv6tSbXeqeLFJ2WWZ2
mA47FhLigJOr+QAPDkwyKWEHrUMNePiXENPSUtXCkRxFbhlp/IMfjWUR7rsH0hoiTqOT6n7hbdRq
z4eA1WQzolWRTJC+nq5vFc1pfDOni4VsrRgYgbrvXapJ/Uefj/BXBJMB+gsqRUdVayFKuaBIbr4R
m/4WCE85px2J+y7lJuXJjnqM7uE0J3t9dGDc03R1srvp/RCo8dStgmx7vHcmcO9bRsaps4NvwuuX
0JE+twoNqmEdyFoaOdBqTVWWgMTCf3UtvJnqXKTVQ07WqHwXS5gmOU9NX7YMK+Rw9pgRY5fQoAWX
SDwPoQC6PzinjqCKU3DpssObM8Apj8InbBzDZPmpDzFmncnXwxIl34063I4gTLt4uBBM+uJeFKXN
kYmK6TcdLE07visIA4skCuccM7AGRO0L0ClKY3ShH58C0g+5hg2vaj5BAjGrnzLrrUQeD+n+muyg
Ww0HO/DsCyeY7hTn336K84i8+U6XR19yRFgGh0ZoQfmYrY0kwGO/hOU8gd/uJF8pwb13y2L5Vu8j
IrPmdEfgIO4DFnfMtnOsFP4uUFn3FVlgC2MYtCWQX/+hpPu2AWR+e383SKb+teDTFGT7eesT+9vj
Lv8BzHxtO+IPpSxcn2KmERy36tUURr8TSBCygK4ru4nEyGbRLbhyZJM6GKziLzXO3h9rIt/X4Aj5
D2kHXDszOmeHhHRqyehpIDbia9ZVlJ5r2Bb1uEqThwI5CcClhGS3ojNAoxoAJRbcwPs9YdMaa1CG
id2H/hyT3pY1SrE/HWDCNJC/SY/TCBNTbNibD0VE+EbziAoHhZ06wt7dzgl9KeZd1qC76eHKKmli
aopcbCcwB/19m9eQc2FJEGvkYnlTpdrwWmSF4ircQHytRi6JDrgTI4MpU7RKicRCRjpXBKZpjtXm
t1GwThNsxHOcxqjFi8HH9CzqbcZ9/JRbRaVjPnRmokZZpqWiyFG6URVubcLZ6dqvNspf+U+KZ4hq
JQyNtwDyuKh5dABre8wp5nl3yBkItOETqBfVPKKfmZNMvZw1sGQvBGydRpuN+8ELs8o+4uhejWlD
U6f8UdvBkjOXAjEd8CrFUpLqD+6tzINt6J928RjsmLQu458hs7HV4LiOpu3x3qcf2ovo4EI+p9L9
EyLR1PgzJjIOUxuodeChx8cSrE7bqA1vZF0GhyGn9+gx85+ZEffXcjb4HyN/7huB8i+on+FyQLDa
5cijw3jHcXDlRu9vUjBJiX5Zuc175HRYpJUo9cfBaoHcJv0hFAERTtYu3T7c6vJ72ZWZl3t0fFLW
uE+qotGxhAbIQnjVu7jjuFhzGALP6ivEbq+C+SsDnMFH5gSMwsj7TwRm8OcrNnKqLYhiGpNaPxK7
y60EVCVqqF03hE3ZwyQHVG6QI230GYsEPzMeXXvPQanmYiPCCrNBJ/D1BVB54PBPiFOkHJ7oWgNx
0iuBPG18FqPYOkepVxwaQSeTckt3DW9vtRaY/hWgSB6XcnmBPCZqdYSSpPSo2PMIDb50hFSPcRwy
FXM1ItZVo0heVE+AgI5HCXLH1KbvRgN81Zky/ezvP4S5GJWbFtg4YVs5gOfEd21oc698X4Z4Mfav
dlDLJFBrxEWCZXEUEkbET//MHCwgb3wKpiMYkAKqDD31INakQVOTUM4/7+xebbTHKmjefk3rtFOU
xJItYMiHJAI/MUIgXoTsTVK2U52WjskDiYIWaJE51fO+5LLqCMDS+X/gvzPDeVhPFnrHEZhmkK4+
57eW4hikkcbL79+QWN4rcr/6/OYjGACaVTqa4WuU3PhNZMmoP9Vr9R44axhOgbWwtkuvbVYZuiMx
kcbMmiLjBTVFWE3wQo0qOQo3RZSWZ6B9ZSRrpTcpoKKVl6SI5h70Vdk3py0t9O8f695lkDFlebfH
o/a9kuQtSKBhAf9+Bj2FdC/5f22+L7CXdEhvNXBiaDS6DeZCh4YOF1JCLD5BHEPBuZSCNy5xxCQw
kaDtSxxUggCvnmLI/2r2XY3YSgKR40iIOxMaSXjym3unMMcYXCey3aPugbyVCcQu0ubuGPZaspPz
GcUmZ6QKaSBYlLZ48t0G+yaufMtsvXe/BCEmGJDW84vpzEjCDSaZ/JK2uRfBomZb5ahXHYaGpNFY
DYHoG9x4rWwYRnUeV38p+P+82xq9xC1cg+ZfGC7tgBEhJAE7GF/4F8o0dOmQeelVOHodLNca+nPT
GyK/Tf5X23SYTV08LMKOyTTQ8opEzDfLXxIZgEJqug8vRBuVxCRzTrPDU6YNSagUNO62DZFjpMLQ
DLcEfkBEeP6O+iJcZOXNApkMPoVPrtqlLdwnwbQY9yUCpnF71v4X75JJ3qYoIOqhlvAWHKlG8Bvs
UwPhp0lLEuFakBE7dxqdneuhtswLXFKoR4bFVqq3XuCv/TtXQhA3cBXtSf1ipchlh7PwLbpMs3yo
C+PZmKVjrif21Ctd19wBzgA/rV7Ng5b+fioEnWNgdxrkQKx+oXygmI+VU3i0SiHDruQs7OMv3jXX
bGryWthDQ1UtKfpYjJ4w59E6YevBmW1d50x9l2iHSR0uPstwLYUbrvHqplcmRfgppXgXisCJR/oI
r4zi4lc117IMjDMRiuopPyiE/6Zq7xjWtehWCY08YdfzqCpBP0LrR3O0/+8RA3BD0LDcHbeEEVa/
GWwp6jP6JUM38saxcZraIMms3fs4oL0P+KP3N0lRlk0uY8rwbUPa0VkvbYbqVc4dbDSqWx2F9EqS
KdJMTyUHNDenUTPoBjPYv1XPZKfd94dgfecCK/6CTbbgLXD9Vw57YybjNae0JkNuW9NqZIOo3wAq
LqnUMx0+m34LjK8iRNhG7x0YlgTRSdMVvyGCwZFbz/MRdim3Y/4gePCCuzMg7eQm+poX+Sfm+AVs
089pzxx3U6dfFc/KWvux5bxmnzgRtIeSxzDXGxPwz0BFRtNwd0bNnu3Jopr4jY+RTOWZ+GsM9qfE
jW++97VrEh7UEV3JWHjOIW52v9vxnm96smJwBBEO6AY2R/UdTQJ+Ji9HoT6OKmwWl8W8fOJwQuKT
EdUcYtmZH2QqEfP5Gf8l5AaVhYT0eW6buwj0EYVKBdqJYiqEDZ+FNIXnm4xq0hW7qE4PNbQoe20E
unAakRXr8Dgmqh0Yv2YLfaskjAVr8uKNQF3KH7zXjDCwxQezQRtzB/1Ly3sFAtaBaIttHWOqUSYK
z86lpPSDAdojVrBVmUDIYZZ6gMstkIDV5OfLys/NcScHUpQURHW9HbJvOXjqhOnYj8U+hkQdor8b
rOyOD+BUBYA+oqHg5u70l3YQYvpIOraPeTJL9QwPSseg66l1/SUUbkKj6dcx3PVxhQbfpmY7HpxR
2Bd+1VOA2hjuIK1OihHipYqHHirLjn8cYEO6Xlz2rmr3yFloBuqWPqyAo7aIAydsXqUfjahM4POy
3jYd19ishyIZsOJkG1LVk23ZBz1Ld69Ju/LJzGWXCi+NBPJ7K7l5ysliHemw3LcALG7lqicE1yjF
jNFDSyOohERWYzBvngnkyX/4QUFsCEwKHcbEwwJsPKFT61EaDCbQllOHxQ9yeYoj6A3AAPiGW2f9
WdEOn7C2UYnA+jHDp635ax/6XZrkaU08ss3UvGrhoysAnigLJlhaHYlvskS3qlYM5+/SumO+B15z
lrgxNfozFzP/B2A+eEtiAJa7mAvK7vvbggd09ddqikYF95kjrpF00LlpHUOGm4bvoFZkHoq/8VfC
KliugJ27s7M/QypUzmqLxYGP4jba1qwQK679pBqTSHV6Ggl1Mg/wKVc9AuGXW4naR71/HrujrK/I
9MoS4yginjSkbMuMkqlJP0eKNxmUq4+bkI7cTCKU9qL80RwyJL4mtJKJa90NAnF0SB89c0XltYMi
tCZvvEzCnxJKt/wHjwh0L2rGEodqHJSDLpW5/JcZvkiy6tSiDUsPJt4e7FRGMln7l0C850zNtroB
P4VX87WRJwgDaKESVArphSdt91d4Ar+i+hQW2Lh6bcaP6XPavgq+LlK48qGbyfAVoxDNc8V7Qy8V
UUduGvPcz8cwWHJqKVrgDB371kpXk62kiNOUz6SOAgPgjA2ClaTqUuh7CoRxw+Nu7WAigX/n1NbY
YxG+3ZKCBhIlXRcRlIa//DlvNgaYNhy5F36aG4vbzmLucDwhOgbEM9S5rDYgYKsXusOyCJbSjJmx
khIik1CFjXZNv8/NfD5f2dFo7n9Wu7ansa+oc5mgMCd+ArRYu5QXGhX3ZFIFk5u7M7dRhO686MWl
Baclka3S+/5acw6PsQ32NK+Z/WHjUclGt+QBp/noqEaqHqHkPbsaDvb8i+dMN8l/4OZ3U7bNZQkh
e/Z/m8hzQX+tENq7HcZLGEg/CpZZALZazr/UTTFaiW7wVO/JMxwUhaUfzt28f7f3FL9im2jIBAJf
FhpnoSoeT046I3/e7wCSnpzojPZsNbpBfMKnEZ/Y6hygZZeQhTC+gasdrUOJbUC9ZV0gdGH7/IgH
kRrDDQSnHNntJw0XeARxmA8WElUtqByLWQAQasg4Ppt4OaMjr0NbLtUcvxiwniuULb2eyamZHarX
sp42zVIr4GKa9GUOL76pu9Bx6vVW5PpG+QnftdIBdgp5OAf1//Oy1y14s8kOiS/DaviOPEAlw70s
WeYxeP7hXM6foFme0QN0T3yMYBHqYlfuPKGWv8m2Cu5uj93rHVXnpW9JL7pf8ZHwlvevcgjF/E10
5wzAph8LNuwcTUwFiUOI5tQg/QX3Ci/mPEYe6VODxQRhkyzrq5GZfsfUGNtmMIX43ZZ/O+vuSdO9
a/6/AuBAzJJNY7t/38G/Q1ihXDpTzS1zbowccWO1/kPXLtbhgbSKeIPqSdBLen7dvGxZJZg4Cxv1
vIxcEixbhBScGJewF7RHQOqXYD7HLzd/BwsfXomxHNLJrNjKTtTnK5yxZppQm6pnI2UFs9AtCjrx
GqNg/l+0KqxtGMc5GyR6H3kQ3qxm/zgiJVJaLb9lROpFpQbJtgwQzTNf2DvqkvCV2U9uixTQEy+B
Q8ucyn5ZqCzW8vsSHQ5ZuL1SbFHvGOWB4FwfwukgVup3mLypCRqWjMpVeh5PaSvWHJ4JQIhJFSl1
Tbual/scn1cC8RWwEsLYVY4zHcWa246ytZHuJ9Fvj3zJ9CwCr+9EgmSTWp0ni3tI0eU53tDDDYyR
hQNq3SL3HT9F5UPlZJI7HuIg2P4KiKRjTQM03dpTl+V1dYUY0j/782S7nnPBj2x7NK2YRf3EvH6X
gAtyHdZCcOeHbt9Gap99fYihUuAtaKHO/FCJej+ylDUztEFRPEL5xWbWIfx78jIsVKTFPSHEl7Ei
g5oQGt2edhfNqHWw5ihAHTV5o+YfDTegmCMgNiGz72UPPBbY5kXsTrMNQuCeXfGdfCoV6DUQx5w8
GFmJVP5YmCESVF8fgspTMI/k4wxHPwMd5yKXPPgU9Wtaco2SEXrrVxMuMF1F1i1GyiY9YAXrtgGm
s718WUOc5VtVL5+zrtRsrTBOfFKrebeXhTGm0aDeal69sXGIkDCNxTuxOg0GyO7krzxXUTrmWrdd
zyjWVL/uU1U6MnbvZpo4uuXzMNswqPSuQ0ZMGtZWHDYWLxb2TYoRUsPoqJijjMcz6SiI/B6MZIK4
cyBPR6Ebk9ijbGiwCh5hW0bXlCy3XaeHUbfZCDfSns/SMT97ogMc9j0aPJpN7sdHWthRtk/n1qb0
+p/d5VV9BenibsCoo/x+cTJnR+gVCxugtSCPwQbitvcfxUmivJSOGmN2harh/+btW6aQSeHhkZlA
jM3OhKnHabbZkzXKGAX3kX57tEZuvVIi913Hhv4GVSrVD2dsfuMm3RDgwwj5nyHR8X5iOTwXdd/w
Xfb0ILasBSw+TpR+cacDZhKDDpUhPu8sQym6R/7uBzcWnNjXCsXNZTzYU6EVJFR4At0+LKAIg6Ea
kogacPq9nKoWyWqicCSzYsw2w4pzV9YnNxpNJaAN/DGWERjPd3dsWBGAGOhPMA2QrJDypfRgVilI
+KUZimGMlvYsrWfggw3O0cncSSX6jIU8NwC4v3XX7ARRF7nPKSNpDrto5saBpvMHGa0h7TpuDHZc
A79qGwx4EbTe5CNoeWxa+1FPSy41YyZP7UQH2ynsTRrmFH5kf8Z+AdQ724Y6II7Wv/m1aq9EyuQ6
/WTeu3AXz3zEIO2lcbX1z5nQrHLJbdmUxdt6vrIg1dlsH4CRUIKpXdQBWSxg+e1in3DrmAct7TiP
hL18YLPfGHe1Ou2YQA+8ZNBdzHqvqAerM7daqYgVNGK+WaPoq8zb8PYPpJG4KezSRLPcc+zNmRxs
6/+YqzyyYngUUuf5n9gTz4z4V5tlJb6dVytz62amNzIePltI1BpNAObm5/qW6/5hJWMjRVHBPiNh
0g7m1wsxhcSzTtwTQ4W7GeUjZpSH6ARhehHh5hSE2kQug7CwCyNTRJ+YWOqrUHbjEbMjSFD3Jbjx
VbalE88cEZzHz5HwpFufisuDRhf5ovzcwGqcnptx3ClGExulqULyMVX2TQWcCMCipoMaUNccWFfk
1BN1ZabX5GwMl1UnLcQWMEC/1yYh5OphMUe54WmNHBMlT85nmXVkjYhmkvfnF2tPxaLRaxDQq3YF
RzF/Iwl21dBBMR6IUIjsjNBOam14VS+GGc92oSIQ9urVCPx8h0vf5b9FPccClNx5NYDkdU4jSdwr
t5WmRq1N+A3qNklyeXiiiq+2l+6yJ+pCiSB9Cat6M9Ry6ymVUPGTCnARB8xcou1lN8+h9Nb0Lq6L
9FFVKMtq/7kRcXuXOCzALR7Jw+OoLteGGltJ0tg8tfI0QyEWLG2BNXjtrCBkLCFYaDHZvtxzQoh4
4TBT4WD0oAnwV0RPV3JqcaQY/IiGVR1ACm3qQlZssVCrVEq5RMB1dxkT44Mphi9/sHMFsxBWaBbR
T7BE3HaU3iu86I/zso6k3qogAbYIgo4+q9OL9EIpIe44X0edVnb9kaIi4BpZWKyQFnDzPwurktBV
pVJsQoOzeE+jdKHpPgnNF6goi/S8gDbmm4MskrZQAUwR7kn5+QK/1wwaTw9Egd6Z9jmCFH42n3nr
eBmFzLoDrStvj/94zcTFIq6ia4o94g5cI5pkRVB4ZIavTxBDvsh9JLSAp9AOkmTox1u0+YBj1Nzy
UG3ClPc1o8CzzoAejkn3dBkfWlU1mUaI51COgdA3aEAUnfuN3WOLSaZ3wm44lFEMHiNrmAa5Z9H6
c7yKO0dQwM+7gDgk82cvGA86vcTCQMt/DU8qKVdbcArGw/fJTU7P8SDINZfFywifpSkw7Zhz4C/8
8TuPNFDY395DGeFVLkG1hALVeQ9Vp6ZKwMDHxbNic7iCEnNf4OpmVlChjXgZybmOtyot6F0GMoeF
z/R97zXaQw68lXLqVPOS0WNbmzg296tFS9Y16Ig/aVfAHonQQ+2/ZjIsSuMsiz+kxIuKaXHd7EZi
VpQxf4+WKOhLWk+cHC62fb6+6kEbGJfx+xqH93K2sVZbI8YU4OUZlyeWx8rCkGvn3cF5gLUXrvNO
8FD+UhICojnFcBKnBJdB0QVBy0MQgwFsrRzSsZz7Q8AMarZGqUZ8anYmwADRrdZ/cfAxKwSv6AHr
6wFkOzDjnLUdjdS9aFN77OBcyf91Fm6sLlCtX97Y1DN/RRuczOmqpcuTt1jxvrBD4DlUGA+GvKHe
mPHsArPyfWUkZdQ+WUjZhlh78pC+ZRvT9DNANwNGgHvGBOz0J/VQY8ieqOyer/xFzIs4UVZeBJcv
Lk0XZKdEQsHhzl50Bdy3fPEj8DKCJih4yWG69lpOLqmk4eQgJSwQTv9xb6pRGJeSqxWcXwcJ8sz3
cl2gVocR1nUXAA8NbkHyC0jouTiatRDOwxZApYMvaSZ2dt+1vXPEE8hbLM7HPq58dz28y5IQzf+C
2NB7AI8sgCVpFWnmnx8q/UtUCnwRMkqdvAM1bN368/k75WFnfX7qw8/XjUNilPQOM1DRdavoqvkR
1OLJcJCOQAzy6iE9JJEVX2oMHuZk+i5U+RxyblWjl72PzUnJ22IghUHVFuFR6qoPOFno2lDAl+Og
n9wWZToPFBZfcFLKCq9lfy2ZdU1yVeujNfVlzdFP62Lu7tOhaXEMiwllYzSxEvtFmxZ2M1rXyJvz
qsZGb30ZUz3eOTSUwB9YBzlAVmwcMEehpYVLOAT9G9da396m1peBGiGHh2RwUP2Eh+vi6ZGGH2rh
LQrmiOGoxcP9MMwn2+sMUrhXLNU+QVtHN9MBgecMVOSBVoXWNcubIiuP0DIxyi6tXQ602GEzGuVS
r6IrYv9bX1JQJ4WrgGLGm+ckgevVc9lqDHzL39wBOJaHRsjiu+eIMAGTBArHuUKjhu57BJZN0JJB
p5PfBI2BtXN+nYhvGov/n8f49xVcmu7w0EjzyX3Md473FAnlMsUSMGNFaxj0RFl/pya8J7klfIIZ
4ZIx+69Mz/NRqV28xIV+mbob1kwAxUuI1zbt83oo5kTxPSqIzutmJdmzcf4SI6TUfJlfmpmuM/+t
kdC/V8L3NFhn7CV98z0/AjEx/Xi/yUfwsjYzuM8UBn1lAZrkAZZPRsywBoCvlU92PbAXHVCyTaVA
erVKbxvIN2JXOHwuWbN/jNpeFCZ5K66XuFIQOEisJBybRMo8ofXiRhmU4zzfIHmHWJYXjQGKXszD
gyx09Emty/MSqn2rBmNbcSWmo1V02kY0Dj22Lq4nxI1e1zROS70VABR/8IIboDkyCoqaHfFp1/c+
Du0sT+Dyk3YOONryG2yu1yQOK6jmjWXrqRMS4zBYSGpKtDeD1uDYwfeTOfjN0HZC7l/il/tzxu02
aDFRteNKLLChABVQGsCMi6Rw5a2+ZmBpI1noC/FRYFm08ffwGTEyo1ux7iUsPnGhSWW/IZ1FYTzc
Igg1FqwnBNT4XnAGV8YJ+3B0PAT1GQZCEB374u7WpF71lLCixxs9hxW0hpQUa+vy18rVOQELjXf5
sE0+eEWxt8Trm2GZQdP/G3PX8Kz5Hv1/kSM+RmdLxWMpRuF840sHoOW+NFH3fvVaiN4xiA/mcKrj
yfziakvfDY3/2KVEJ9bHBwP2MoR4C7chF4h3Rfh2JaAre/784UHXaS4cfj4cVRkMlGbIIP26ApBT
UgW7sBlpTmfXdvis0ZESj6POqDEaIUaKVTEYY5eQuhHvIBVXAIMqmhs0zcZsVoJVHW4AGJfNd4aH
9U5pfqc5eQpVjog6BPRFnVrSj7pbo/+vyS/lroyL9xXGwnibGwPQolXVKgzxe/tg1nlaoyQwvl2M
iFGqkIRpUV6LyHTllilwHnYVCUpFsjPS054YGw613Cs2k2iya8H3ft6l62toWhEg11jF7P/CSoXB
boZEhchCkP86csoNmNzCqJMgMDddscWZ3C2dOPEfWKOhOLaoEO5aE0gFDLjE8lasxVGnPdCo7otr
dfDj4ns+3Vnah4K/wEuXXcxhVMfXCjmPTqmgaekqZJPeSof5FQeY5JwoSGY798YniTSPvWm0drCR
lKFj9wQlxa0GrHpjViem9sNnm5GopqC+HXcUS8n0HM2L3AFimar8s9DPYyr9nOQ6Bumv1kU1F3KT
Ader+wQwPMDJAt2q5EDFi3IR8TPalxBdRXk+Dwpt69ygpmpHAkb0o+ge2rS0xtcxJAISuVRVUaqm
u5zQbpBxHhOGm5KjdTd8wl6V0J1/9udxcE/FK90mXrPVIvHAsp8N1DcVl45rS4FrB7ibDg7OAPfi
3OQMqgKJrbu4D/BosAg8vGyLT6WWBSGS3+jSprW3fYiea7oTLuHjwHOJO6IBLiH7fnWnUuu5cGaU
YRE+xIeAjEsf3rn5JCOVit5+J4ijmjNga7mqz0WdBazIDx0NKZFUCriV7y4madd6XLrEQJxP7FGZ
KSqv/ubfXj0P1/kQ2huirrp38umXE3xJ0Mf/Md7AIimxn6tygo8R3UjEMcI2XBEVkJdyT2rr/U/R
ES3JRTEscNqPmASP9YCTbfaZgf5HMCyWAG5UITSiXAN80v40rDDYgG6OhiR9+Piw0y4DVgFrSoI9
YzqhZAED8GH6Koe5hQxKUGgDo07qxOmC1+NnnGyTaUrTlJAnqVKMCMB7J4WWvcNtMVJdXlqC3KsT
N+tJxzPpMpKTv0LCs3jGm1LaiYT8pZUYWW+h34+Un8a9JPjzEUU0m/LaSm7sSz7alsOJ/XDv5I9K
Xg2t4Skgr8CoEeBDQkrXRIl5bUksrpqWPz4fCi9cFigLTcFtsWc/fgRXztDN5ngIuxzzNkBh/ptA
f3FPnthJZtjZBeyubD4Iu5LZ6tZyBXEDnKxF0Ck6sJVmte3+/umN661c26SS7TRFPoO7bpnzbS0Y
HAwQQ/q2AtC18f4RLG0blfKAvICILR9bzGqZYZQcd90QgtjsUG/bEmnZ90ju3ktPJuNuVooautUF
k5Uvi+rxRMmbhqSrXegRmLGFNZLLm1j7r4aAdf/z3SW1wfzUrYUPL2vHLfVJMmDenyogM22kfrWd
LpqyTpLcvARB2D3pDA1UkyOOPTMuuOuB5DEkEnp/pfxaftzaSs6B6V7FlzIcss35TM0+cmF864Wv
qjEOIROiilUFGbDbPYyQUcK4ih5AFS3/pCzHnBQ11IUU492vOkuBGCWzRcxZHd+p6pYzOTDO/fzc
H0FRcGPL2TH4ijU82cYmZzPSgGuk75GIhfDKbE6UpkBuOKM+yCXtrp3q7FPrZYgFg6k2AneZ5dLF
GfsCf7gCP5XJrljvFv/vkMTztrDMHH7DnpmxLxAYfcpxyBSHWEEts7PM4Y5HU7Eidm3zD15X2P9D
hwhXlU93z9dwwp1Hocshvgv7FtHBG37HnlrWDdaVoh7yG5c3jUr0dQznVvwJNAIAdtgfq8H3i9ro
r8C75MWCdXp+h1OJOLMod4+NPMhXYZ9qNmqkQc24Hmv00W5wmKeQfzA5lgcDhGyZCvEnsx7pGws/
3AIX1o5ceXVAsipVYzZ8N024sJy2W5kLDefPQL//GI8tKIeOz3Zj/ETf8BsgLqS1qCmxxYglSsUK
U6uUK+EOcLpTkV2T3z4FX/XR7XpKVvWU3bhqDGBJsdBTTmxo0atU51lnspMvGL4m1Lig8tCi2nkm
RJDlbv6qsctizFBhm+HltE4Xu7glkgKNfPd8kz90McuWejsSX3zKwjJbme7GV+48PdBbl26pVRco
9bmAKaep0RJdFPq1KhlJJj7fZpTn213xu98tptivQ9zoMXgJqlJ36Y0uW4h2hbnMQgnjkbc7DLoA
sTVSA5C4TSd+XGRCpySk+OmmLkhRrcnzle1nn06M0SxhZ+wuReyFkhDbPgxfmTWNfgWBEIyi+oQT
0JjUg8wqvsrg2AnZVGYN37mK+tfw6zbTgWf3Dkyz6q0CEyFUujpwIkaeScWn+TMN/eqU4vvX2kKT
QKhYt1HDiXr/WHRlLmTOa8EBxvGC0fGvUuPmR2nhRjV74ClLYdizw6u6WTrVZnN1BzX1aM8gYgsV
HbVpv3WCYHTX38BBSG2REfBZZvwH0erpAsyPZsHrOFxP42PZolEQlwA5FESTyIX8MQV7Y6zgzaNe
ecmGxrNq96Ujdpu8ZFZfEbo0NVCxB6YrGUDjyq3wg5OnV9tEr9XIUEw1Mu8JHhk1lvKAzsp2ePOP
Iyt79uKYXbNp0TfAtL5ynkp8kZho6pTfZiumYVXoMlmKvZvi1d9vT21K+4Wg/birR0AJEgjEKQe6
N5eNNahexlUfTKkZSdKoq8TBjaPvl+IA/uZF520eJUpnP0r/nRBHNfoYG87heWyQGm2o0okQzU3t
1goKYDzxvEStsl5Qh8NCs0AVAgnmJUZBhX0mCFhQNNBkjB1KUviF6k5dxrXuMBsfvzfp6juuy8ma
jADamPfhWWeMZKB7Dp+DJzhH0yKxeMHy/OaCCJuMSHIxCgIPgsiVM9ZiRmwC5i2sUG/Osx+eyuDa
BHEjzP0sMp2Qwjj5C6FopX3gbPumFs4LdFORibKMke2yU3CDkSnwG6u+tqmHPHvQOvagsU+XSO3R
2Ri2JRbNjHu7BRPeYwraCZDT4tm9x+92cMmunEO1UAD3NKLqIItZStVYMM9UEYW16lqnBHldW/m2
khjkYnvlJ+AFx5/Xp2FPrOTyazJRgTwt2T7JYPno0U8sCxD2OSss3qxr72EnxnTcMHi5yx2iHCq0
bXXnH7M/KzHuUNj38GTp/ZY7cG/x0Hwtlhn8FKLpwV6GwHcDtWzoEjbmeR9v3K/A8ePNCYuKxRUe
glAngf2/eV438oiBkqyXu4lAVUXejM7jHMyfaFuWgx+nVacUPOefBEvE/EDydkkdrNG5/uOMO+cM
/YTh6hM/icplf2qja2OF7OwSeYIzMViioLeTey21NEl8ZjrTj+Cg3aCvHAyCwR4AtECrV4YjPgGZ
u9T1DTW8S7I5fD3Pc5ErVDwx3vYXMSYoTZmSR9RzGm3SMMGf2/3P71agOySL/4A/vLbgO598MRsj
A36cEfi30B0F9HVw4VQJVYpX/HCg9dFZd81rvQsYPXKoagiLYbzCyFrYT4CGDL5m4ERC/4f0U578
mg1AQlHbtFRJ/xfmwtSJSesPexEMgDT+C0AuOfjVWgKDghIzr+wDqiRI5C2/Gzc+T+2IKKuQzoO/
02X7bybtt6TVRHpaNyTHfHwO9HqXt+2S/4IO9bV74P8K1KfgUyCPlKk5b+EySceCSBkKGKz2WbUe
S1xlE0OS8zfEEP65eItWlAqAve0kZXM914n5pRRYVtFvQ5OM/lNwejkyA6iim4iLQs0Bj/KvJ0NQ
xf6kMhFDEi3oBA0mQ9LY4iOUX+pdFGzRNakeIsapTuMjl2OU0X5TYUknqK4SSknAoW8BkKxEKShY
KQ5KnRd7lSvIVBiwgkllQMQkABplERzAcj68SUwovyPT/X4SrlKmGeEWqA3tkkDBgkxooIlVU+Ih
Xrj62mng6sz0a/16aUgrTyFvX+5CjoasPlxRrgm2bPKT7YSw5rKRyOKsWrFPZgYEjhyFa4GZJz1q
UroWYjuH2QkkNRxTkhMZ5RmzxyfOPhjU3jGMvLc6FBkr/gkaHyYJmXwp2xED3FxFehcxjKOF+cco
zjwIlt7dW0WK3WU7TY48xLk9W8t6Rje/AWYyj+xmGOqyLSEtg2k3Wmx83ssoDmYA8Qcq0StQxnlg
y/XXurzmPRpm9omuK1bhLnh4ffhqnqK7pI9tH4BeWOEGCYbYvxCv/CVmLcHOwh6Ad7SZlij+ma78
9mlBOQmjMoxg0GRh2T+JZX0UYwD+cG2GU22hOgWVictlPtWkAsOXzKVUwg3v0OPSWAp1QwGNHVlT
zd+TeDYvI99J7bL0DpTv5zs61L1dbqYq5g4tT8oqMsq3jfeOfOcQ3JIz94fM3+PSnLzjMrn3EizA
DXbm1pjE+m23Fih9W8EiVtzGANado+valwxmwx9D2zEnLeReIYHcMvbYERWQtmi0ZiMr+a07IaZZ
UpPka620cxCsUQvoxB5pRdzd6sMpZ1AXoxp4dKXyFr8ceI9wLyY9HfVnKp1uPzE5s0cmA1z3sdV/
F/VKGbv8f3RoRtj1fBeUcFxM/1sMBaJlH3nD1V+IDqfpgNsbVOyjyZh14RPwIVTVEbHk3Yu1+AG8
K+Ekz1RIhnahHWyCXc0260hOzts8XBsfJUiSDNEbfN43c0iZrw9gB34A9OSWxNC1KNEOESQBpyJJ
GQjnbyYFcn8XxIRIJPTt+7wowvNfGwwneLUTGCJffnPMS2JYSOP872uoz1lYsoXt2KyirlH4JuGV
/Q6aPNZcxyXtzV/vScRpuTYjnzksf81KjBq0EMeUPtWy5hPRkpGlTcpEXJcV5BtCmbEbx04NrRca
XB2CY1FmzTysJry6wXNeWduiWQtTFcCfNF7ueX0oUaigToLCdHFRoy035U2FxatQHiDd2hXnDIM9
bKTYwGx2Wd2D6dOu5nJ/F2nacssZxxUHIo2V/Xs1vbgg3F5c3UgHvlD9cj22ixFdGriRVjr6m+yX
9u1hdZ6YHR0dmgaoqgg5wJYWvHREoNSKMQN2usG0B/YevMl+wD5lG0LfC2S1RjDQFqltAR6mBB1j
gDh2QJp2i0Sk0RFlW29pioj5fhFwyt3WMWuhB13TyUXwW0lcYhjdo6REAsFUngcpw3roogPVgcrV
t136GxlYeQWV1LBtdzpn8KR5VZwGs4duI0S0kAuF4Y3c0Si/IQKBgeinlqvHou/pjPKt+jbODKJp
Bi0jAx+LR27FOg+ZUp6F6ReWJJgjnk8zG06jAnYZHOga2rSimCV7F64WynO85VJHZ4Mn7onX34fm
uDeoxOs5IRIsh4K4HX2zTkq0bSq8iiO0+3XsNC/qGjoO7KreYFR5oVEmnvczUpqT9fZiiCGPamSC
1r67AVkQxHEP6nR+MxUzaLLF4CjpHhC2mIE/RdtRAd7lZlNdgkZJXjI/9/bJNp8XKP7TbYwkwfa2
3qzITFMErF6kD9pLSuz29u2RhYXWha8c/pJ6cUyGMkQHSTts35NWXoBiEd7Mqj3Ktk3xo3jG9WFE
uJAZc5ZHyu15XABh/3LcMkmYE5risy++q6w/6hBGgkx4rXtM+BZ8B1AYzQbZrVyTRmxQ2qKr9di/
uHkGEmbZPT62nhmq2AdOLZC1D8QPFdnisIkaaLlxJRzVPWcbvFX+bFRoqznKiJr/SxLMOnw3fu/c
2pixQw1GmAOVmuRhsCiVd+2vJetVSZa+YNQkeM65tJ94op1mZq2rZJ3NeaXSFqP43HGB64U16h+/
Z6w3fmvFWKE02M1Ka6i90mzUbLKx2jy2kDTRHCMW/GL0CWGlb2OfNPGqp+ALO1i1mlFq1AmHVkC6
IEZUu85eLD31x7BTTdbx9qSck+HR5CH2BXy2OJ/Oc06ckk1yzmRD9h1Bmbj1JpzOzd7mhqWfwoK/
4WQ302zxLBPt7U2z9KTQCb8chtBZeJ6paclHlRvc9AWzKj4UIlwA0LybRvEWYLLEbyotcIcIMd52
tKqT4c8qt0xxNSrcCZIbj3Ai/Sbepe8HepDN9/SDdwI1HoNmz6rhzHmLB/v+c3et2LrkaAHxzJjV
rpA+h3v3r1YmgXpY48rbK6SrnnFWrOJXQItBWZmJsmfsKWI7ZQMIcNwixxTaHY8c48Xwp+FiuWaJ
MO4VnuGGCRGKwLqTFcwR+/UlyzALfW2oje2Ez3K3S4YFnbwX6GFDxETzpovjt/yl0XWqO9zR9LVR
Nj5ScbB6wJMW8fl6Yli30OtQ6K0Tj9DRE3zyicEiWJzHYdmo8qHqH74ZGMcmT1efR2RXh9hXVO6y
oMwlpL0jt6yPaLAeJbsznEVPgjW4gLKh5zqPO1Ew7v1muYSsrcil1hkPQHeJ2hy4rsbhc6KJVp3f
qgHPxZ0xL7hTveLc6hlrxbP1m4i9IUExvn1NdWNOHKcHyYA0ZkSJofvneAyKYTuQky4ClV/7fV/I
i0i54GWKjuepuj/JAG6ZNnX1ijC9cmh1dDYwrewDKqEGru/mvq+hVYvPJYlW/XLceTZlEOGQwLUD
e/L+ix0zSgfNNiFSxHc/7SF2BFROPZlOLMCpJ8prnNFU2IQZJuv2kfib+P6CkjqS7eB5zWAI6Sr5
pENs+qoxxw6hZ0qkDEAJE9f8KYVPzccZE/Z/b1mLOcrDqZnWHWH0ZhgHkmbkFUGRLgrwJ8MAhpPS
4I7uqm+6atFcq8/Fx3GLFw/ps1+v/irObWXjYvaivsj3vLly1dvaicqLFJk9LmVmYIGXPwQ6djpg
qTLzJqSiI1uGIo3QNNI2Wot5tyiKXfx15piQ47lXVddJMI2GppYYtaH6IyDtWhu3O6KXM9uQc58g
2O+mimBzGOexMSGemmYaCE4+Rfe91DwfIXSqTTYmVSf0zMP9TnR1vBPFUUaYIIKU0sRUL6tuhxS5
0GjHEDBlyFKPB+8Y0EqJowV5YygJYobSSJ2NNLifxv17wfAsdQyJt6W9RBbRhk7LOvTBoaydo1hc
aS1kTK/u24k1Mz3yHNcmq7JKFLBCToIswz8sUOty/tZwFE3HJTqlUzRnYm+g9Gg8aFdQMdRC7qV8
mmM3N2XZhxD3ibqSiNjqQjZY0ACm0MMCm/SbaAQfUb2QoCmkBP0AI5ssMW4YdrE6cMVCls7ffrDe
qdDUk3yb4wf0eZaZaOufSeR97OTl0eyL0e8CI7nPLXHcCBRtqqACL/C2Gl7E8QU07+1y2lwoukcN
H2UfiwNv6/83FLdnKGo0yY6vybEC4H9wdVWOZHz249yhgj0UXzQ8hO+7umP38Bam7lObxRBMX16+
BUpBL74eheVTwOfMMDmqDd+baNFbjPo7vh6NAkXO1mLc9OxC2fZMLD2k1amfrR654qKu1BU/44Lz
BCAGxUgF/wZBFfRzeYxafjCpiYOmv1E6+gU6dCsKPu5HdecekQHMdBQywsvLhpvM4KxvtS8FVsux
zyzhzsLIRaCzp7PTrB+AN3yj1qeJ9MBM3uDLBDo7/5vWxf8dZvVwfSTl96RFNbaJtDPTjVD6+Vis
KMsun8MMkAj7q5sgoltZL3LDcRsVJjmrELIO51G83H9veikTbru/HrArkwlHMIGyTYAY0QxHQLIV
eXt0BOm/t27zDuQnus9hhRaF50MGyIeIMsNM+fDeZ4IwRjjj1AEoJMfVLGUmSuLLJMcdA2UMM5lo
NQ16jS2YeHK3mrsPnLJoe2ABnYQawnFEKuNzDuJXRWHiOlSIAeZkYYEf002CYQX5oTgTZlH4ocau
ltVcLuRczUaHhp/tInMllBN9mNi8fKztZsWd9EHTdW6n4TGMm5yhMFuUNpTAAK656ca3eNxA9p+y
HxWjpSaep32+5sIHlBeLIy6G0dDrBHEZ7HLdVNFmjxOojjurbD1tAzcpRHZU3bTwRpq4QHEUwl3Z
V40GIz0/qRJAil6Njs6r/JdUD81SO6DVJ7NlZAt9NaE8rTYxXYz+YmEQQr7ywuAtNHRtsFlfX3BH
1tyaQ89s3OMBZ0BVc47Yct45tcPFYXtfuweR+fErpCJAlF5rf5wF5TGhUNF6+G466miclcabZQmH
QJfau9zWsdXZqkgfmp0uL65hENml8hlQvkMhFy0FxEGitXBEfURX1QqmnDVrVKJA9FwppmOtmced
alC0p1m17VNsZ9nyG0drdqJahu3W5PibR+CjXnBEgrBSyOh0XuGBMme7M3q3WOlYwRMMwwAyEMjV
D1ajSueXM6XGCVehVDnHTApXbRWio03H/YMoqbj2YXin+xIAoHjYYFXEntNRjC0zKfu0QNjt3uag
zBzmHRF0cO+le3JSI5ACg942yv/ItRwpmCERgudzEnAALcDi3U9zSjuIvsoaSC8HOLVFhbyHHHaI
Eaw1Tt7cGk+Z+te6FND9oWarHFLiythfcslh6gf9WpMzfm1YXxkQjh9zUq+prTKQO9OGT92JPb66
MPuot1rx1nMxb4f0cqjdM6KuBQAEjV2N7/KCQLC1DTBvkUnhWRKM2nvZ4tOd3SM4Pgu/7dmp8FZf
Mpa+LG/t33AkPLdBfCzSnK5MynxK+MTOuKUNVkwWdFhKp8awFOosIAa1PGkjOUT9DbfEyHmMSyiX
yaY9gaI9IuZafwbaSYy9Mc9NJez0fnpsTVVlaBOdq86qyyW3k1NRis5QQknnLw/Dz/t4wW1+UNmE
AhuamzMxpOFXMebaVyYd5gKrtgPeyXqLCiJjnMo1jp3DrxJ9vbTmCuOy12DKoCcr4zymfghXuNss
wk10yWbtx19JBeTyOHCx+DTzH48NzWrCHkCWyw9BfGG8RYM5ke3MLCvrP3HpfkQLlsu1ANbY+29Z
B0BjLipoGdAq+1Pu81A6s2Vk6IMFMbDdRkxQpTVNX/nWyN9FvkDVoVGzmvpgt4V8Yzc50o9vwL2c
g+TlzuHwBkVZhizTSmIIR9FQ2BWmT4hKn6BuFvjbMfx0ExgkXC974dFUU71PzjjDWiJhoj7Sg/P8
HIVVe+tWfCLaFK/Dm9gbbh7LbJxB8rQfvqAy1lC7lyhVf6SN3wHkvK9MdjzUq91JKmN40TDsikFW
XbHK4G8Y+Vo6KvIXjBV0pFazPtxAecY+1KnO1LkcXLbh9TcGrpDxKiTDcKx6DcmFffrBnwOwaTHI
3GTo406FEK9hScKPmbNnFMrPrK456DWtj6JFdAA1Urqh7ARr2uZ+i4UnnaMfkjhTzXX/+GMmqFeK
qTw9odb4Sof259EXaqnJFIAOi8CKFozLJTrJhiiy2/rJBzhHEONuEcbPOglvDdL4/XTwmp04iMWM
KnzilFQMxGkV8ZtlHYqL++5DUKCbVIbM0KBFbBELiBYICjgYpwJvoWzfKf5XxNAxpcV5yDdCa8Re
DQPPOeXJaS3zGjrapy9UESep1YEsfqm/bZeWXy1ua7CC7rDgC90vMkTodZ6iiH3BcvdtXnHZ+LR2
zC0N1p0fmKrmBiD9Qh0wT0Du5IMoncXGMHP4/YX1JQIDTn7TwiYonnsKF6PBI21Kxc98nawMKRKA
2O7pBjv3Pfy6AIglkBHj5VYhf95NieF1di1qnwQqeBZ85UElV8CIWkLafEJHQqa3Zg+DZyOb1Lmv
yFO0j6Np4qqzAnd1sbpih12MkJteh/DOMVntuey0ZSXcucgW7TyEAMjl3rr/acNZAu9qB44B2t4o
FvchIRxldPCJGMjTff6c8pXA46J2WwaI09d/cMSTde4Xoc2hEFyOFn864UxT1IECtXMq02MFtswV
0eT5mOKdf3UbUuw6KHu4Op/g6se8FRB5sj1skojtHKaajRG+jhBcoeAQJsjX6dQ1VhTat4p7aZAy
C7eE8hIlG7O6H4umEKtKNZ5SMbb8tdOpAWIwct9+QvAT+tuSThwrIJMQYJii10xfH+p5lOuqLrIv
5wEdIRV8L7Nx4GryC1BnPw9HalMb+8Z10iF72yhmSVIDt4MnzdJICH/a0aoLmEATjpFKjh9gB9+Y
VyIDqPZWql1O6t2X6DHYrazdywtqASjOgybziAxiQ9J3dKSEdenwsmziZRHmVXhDwt+2OLR77E1y
6W2rBSjsX4FMrtHgf2BOluV8KGajH84nG3fxicJNEkpz3RHCrGtDdThn94QY5VA6p5VLQrr/3BaY
DlnArr5Ou2enElpd7lN3Oul2Gp2WFAWsahUTHFHED7gVZ3yIFwKrw8ZsdgqosiI92PbRZgiVeL9z
rZ47si+BX3fTmGgg1ubv9b7VgM3j14Bt3s7L6u7niHFhvQIm9EvYBoJjcvmAgh0J3i3jfqQvfgcf
1136xpeY7qE+xmgkOd0pAayN9smr8PNs2tXCIBWSyECxIMkceNfU7v6wHNBbixJDqnmeCcZJarTB
p4qH+St6R1Ni2k754VGFBSZvlOfmMwa2ve9ux9hPQ5RRm9FMHuWrEqCQrkOyRUMHFoDOZTq2jVWc
tBzp6FFqlKMzw2UyBCoH/3Q9PTgDqnZA1dr9IQZ1H80CQGvJAjQGp/qpOHRremT7WhRasio48J1a
vv+UW0GIB9NT7ZglVhqEqFonq8FGNl+8Rir7N2AbRrEC+T4193+hkAAM2cZxHjV5ZCGpG6dtbeg3
7sI3jtP0hh9GRCCi3fq7r/4OK3WH5tHW/tdpIMG+EDYYFSPGVCDBXlN6JMcxlLiaIurld7trqFvr
2MaX58rLM2kmMWHElFQs0RJ7DCocVcsVmvbi/iC4zSLV2I8N0SP6w8RCxKh8B5DPX+JF2d7fA68x
dl2wEKdsG/fbKkZ+ufcXA55aH4Yjkzu3lZDuA5pQVkSbcjYiB2UshciPbePbFRq7nyPTzm9nsXSi
4pMFCIcj0vhWfWDeX2rqXFjVOrPJvMT1zLQx3w2sC0s8Sp7YbWDefZbM6N+aWL1Z/isXbBDGgiVn
XyzSBz/ze77XoVNRIrGsRr1nmHBPmU4dg9yfua3LSdAVxnqE8U55f42gISTFXbkAVCVQMXbDlzT4
R5hWbFOUHgNywd6QmBSIVFElGG1uFKBwf9J6EMseJwcR3Hvgc2IWSc/Ew21pHCofI2bAnlFDiQ2G
mgw81BHJMBvvyfgLIdbA6f1Ptxcpqb3RGwYPB8lhOvW/p01sHCvzZrOabsONluxJRsfV71UVpcJH
tA5ey08OTYqaQqX0f5YueytEvfovoRirEQyHT4XduFzFfJWkXqpqM6Mw8GP5LsrcJt8qjNMK5+fR
qEx4aTBUDeB6Pu9jPG+BnohAh3LEUjcZG1XENVXE26ahc8LG65YWP1dPcAdmtrBRj5oThHabuVzm
WeHmmRdq4KzdkmMYFliHkHqyzXXGpJ+uzgevotkXoTZ/5SuP2FxOQ3y2KqxIny/zdZBoKHCPdhTn
tcG/RiFnc5wmn780D8vNh3jevZdfpsfHjkHeNNxupZrpujXHiTWI/xqSDnN/OA7oZqJaoSZhbgqa
vJZYwUmYIDhBWSVIwv09efmD+HDPEuERT91nTlRAapdOti2XQwY1PAEu6QZNmf344zgL1Ne93t2G
PSKEoxZq3EFFuOs/gpkE6g4p6G+IrOTpJwHVBAb34JcLIGcc8Gl3Ngduhvfga+jospJXh15Kfes0
SrvdjDAYH31hUEEcSlWk9n7PLmv+PDJ468O3ynG1Iq+9eICMgOWLzMhl9xo9pYBRAdLupVYuzpB3
h5dl5+CGZJ82nzCv4ELPPDzN9uOabf9nOxI7omu7IhfLZfsaQD0KMn8dTYMbdSaeLTbiL8Teakjg
8rCzVyv04A9M0Cl+MBaEvuXTukLX+WVJgq1qK40j2iJYz1TQdEK8UdFGLiSVdCIjRi9A/w1VB+yt
LK55jCH1KDWUUwjnJbBOLS110uEz3fghvTy0gVrOYpXmN5XU0G9kecRMy72RbdbVvpcdvTp/UPhM
+ZUmJWfNJ5ua6RVp/gvCw4wUjD3P4Y4SgEs53nvYDXcglCCQuj6wL1qjgN98TRw5h0cry+vX64Yd
H8TYSOHOA6FM0guzmIVRbGTrDX+ANY3FnQioHW1fkLcE8653rrp5SlFsHpnu0vMZ9j407Rte98Zr
UECoLztOy/rvlNUeJtjmHYNv7SrEUNJCHM7kZaJMeFDmH6TLU+LCXlncY1iEE9/i9+/DVpWwuZ4B
h3lc1hWAC3BSB28E80yKzm3MMQcP6w1h3H+bkdFHJ54F6db1NEO5rf0etOQCsOHVUQ15b+TRIzxG
iKatWyfn8kUDGeb3tT71JAUweko+pAWg7T+38doW7Py7qWeGz75R8HWq97Mi8oU6hZjKhfK1F7SP
gZEx8MYRCJpuhXFgCnbmv5w7SzsbQayGvkCK/QNz2ohYApuNtkLrlYjbFOnKPOsPxflky3C9gzrf
rUJ+Q9kyKgkBXB/k5m+kJN7axh8v42NWQ3x4iYf8X1ag1sDSWHXnLzU1F6Te5Art0Tae7nvqXw8B
jJwt+Ujm+ap5iL3/dijaoLXGuPJGNiyEz+BYa0tJApPbtAH75YwtS8gsAWa6bMwdyctNLSjLqNUC
hBtwq3S44i9Dkza8OgjVDuJyJUJ+vL6i9GEgBtNpfeE61LERtyk18Y5Ln87wvF0jR1x7arEP5sk5
TArox+YH/22P/ArTHjcOYUU/eNEFS73bIWeuN/X2YarHr/3ZFNPAkN+IcHNhrmK/wAY4Pb9OtcwA
n+mMsXFhPGYIGQJtttwZpMTl38jW+xea/d+S7XH6KMbi8uOmaFkyaKBZ1SAY1vcy0Ji6WVThC5hB
KJhLNhy6R1nmrw16UsmmbFR5yhSd4VPD5M8Gb+WCPkFUbbhngg3QHMgtNFbZm30h4s4KgzWwJ3zW
1LHDyfUb0PvQJr1zvkT2Pml4wzlPhnQTU0F6ujQq948sc3M7B/HvNPzsDbgegYBr6wJSgnNMNvwD
lIspdsr+FLvx227PZqeGzDMo0AIFGe2tlcDW8phzJhwOdnrWXdg7vZGy2/hVzx8gS1U+KdrMW94X
7hDpXOXRWJzuhE4WEFNMWiGhWiLhdRRvFsxYCZkGS9At/YZ3JMARAK7Lr0bwOfz53HqjaWNcnUcH
98Obg1UDWsC/Li04esuJHIU6sNmkM6cIJD3F6MxJpOj74Amkt3Xf+1wvb8j2nzjoDFyhrmfeGE7B
7cJA662YG5zuqLY82MTX2t10fKULMJInnz2Q1C9OEpzan0Gu3+w0ueTVMmWr57xXx7CIPzqtXI2e
wTemgF4pV3mlxZEkqkQLe2aclODGfFsg/TdKONgfoNryVLt9DHxOxH86WanjnvtZlXHbAkP7qCGw
tMMi6CmpJ9ghY998Zn+cpQ748M4JEpz7Bv/t6EhVNIAEC4542MMglDMBk1Ba64RpvWTuYh6SqUwL
ERJAEvVJsD+TJzsgk3MV3IB3TBDmN2a3V7dGlWZ0Une+pm+mz2jZBM74CmX8KpJAI4lW1gkgXAnq
0qGMbKpwxAiJu2a/7i62/pEVcapHJBD+J2oaGJPshsxd1p7P2RwPZ93hH9qZVFi6pG1c2W9NtyyH
EbRbF8iTWbLhxDg8KQQjH341w0O8ioozKz3pmJlNyorBxy7KOi/AOxcesydckCOpPwDNeGA8dPtQ
liRTTeVJ5qEmfEHxHhuVA/BpM/Qjf9QpeOBCxPGFa3AWW+NA1HJjOTKG3lMYWeaRmmAiWsyYnzXH
nK03KeBdfnAoP8eQaWhH3If4vtDx34ir/8husK6H3JA25tmGUZ2eIVbQpBU9ncAdOcH4zeBqgfrS
XlPoETLA06LSfJBHzTwhBz/n6TAfLwV0uXz4Mt6ztva4IlTW/ivnm7AVi9f3nFI54n8Qp6Iwyc7l
2Pgv8S7E79MMod7QGhZ1ZKWwxS4D2eV+LIvA8m80W7qHtwISq7RCDnyt5ITA3FLNUOLLCD/6g3wS
SVSv8Ltkn+98LIIVbTP3GXNw2zN5akeU6P5J1Ki66PeIe1I8ilEopXZVuTGz1EB1F6hgYOE5FtCa
2EYeYo9ddOKgTZZGll+evuP+U0McOE7ibFMHOGMNPqpC8Sv7y/yae755BKKVf/Fzwxr1adP0t2ZW
bqZlcnq7f4Dm/Jm9yoHqKUuFrM0pZM8htVcfWI3SCA8U9aYrAMSygvO+t5ZaQH8QYulTO1BqpkeW
hNuKgf+DEiDAPSTqV9RuPuBRqY8gB0jHc6fZ2AuM+VsLEwLQ590m6JfF2sjTB8WrC/3PuVcVkNo5
s6tQuFgg83JMbU4ZAYg9JjM2sptk+qd0PScTj7aZxEl9KXFw4MyusQNdlmB3+1c9N/092ZQpmBbb
h8K6yz6sTbn0fvHKgs2zWJrWMcohsWLYwZiV7UGa9DR+oNL8b017DPbnqYoyDuan+sA6gN3x0Y71
cskl5B7VNGwDyge3R31Uj+rgPOsXZnSKJ3OezpRn/ZPRudmIIwyJcFlxzb+TTeR32KsKbnqsgPyK
ayEPoImw3oySSj8i5KuWlVl7r1ISOUW8ExBHRhHVzUO4F/h+13Yb4mlCHociz44jw98t+Vfv8166
WbDPWX/dIGEN46nX08D2J5i5Geh52TNWCJVZyKqJyfiPCgHwewyaFZZGJJvBAk9XO9rl8tKStGje
5PrVmsxcH/JmpPBCR+B5CrauADeIcxcqM3IGzjNxDmMMBgT4d7bWvitA7bXSdK0s4G5i4H8e0pZF
IXKIE8N0TG9Ucgx1oQtGpbslZtpVzFXBBdmy02e4DbaM4Z1kXLXKkC4mI9Tdg4mTCoXi4x0eYKnF
I4u9n85d6wnWGBa6WO11+7mKO5AB/WN/jeKWeahVCFHCgMrx4haHNZhbJKnzD4+sAnMHJnq2GHwF
xR1VGobX1uOix5ni3cqEa3yl63dxEjDZwOA6uh2Mk5ixDQiR3lQiSk5dZFjD+Qm0neOuH3z/2iQL
9JP/swwnOdHUe9IkdgkbwvIZ3zQtVxQ0Ks2Sv4kayphGB9an+njfbs4wEt+QH0S+W/icq7AS4AFd
UFFXPzgONKyLYNJwETQIZkEsclPdA2ezlTBU5C4wwE615mcnyq+tNlDBZgrjTltrb5W7JnwT2sYz
0a2SO/JebQ0xXSUQRrkujgQ01gBiSGfh2ksSy4Tgl2Vsji7CKiyskfFX/zL6g9nhloUlLJwLPC4I
t2NMiv3mYK6W0bhJQECOFfN0xiBP54/CCJaH5qFiNLlTK4ixq7JKqecGJnjQ+Kld68sWdGXQHBbF
WeMUtEeUpyjrZcOMqIewbof9pjt4q+V8CUhADdjW2F6+x8F7VbbbPjKIUcMXsHVzBAgojcHjSpkJ
7DwUBrwxu2BncavBlsg7fmsQjpQEIf1CZto3oTSfRYagEg3sOXg9wU47etp3hEMsEv2L6yzmksox
bqlQ7c7rKEO18R4/UJxzxTj8Q/QLVK2UxxMx9+2sHJ7qFuI2afhSpG1vwFGUF3vp1JDqMH7V6A1p
Ax7T/gDttpWJykIm0X+MsCDNpSruGc1G73DF2eBwVfoB2niOZlf69hBlXmOWFiIzWuZCxF0hDp0d
7qFyEkUOgYSdniOnMlxfGt5ZZ/ISjmpoxxBxenT3mXkIgsAzZ6ftq5b8O1pgWQ4MSuK0nBOxjgoz
eX74H2Sl8F5Y3MONHVlZLg5l/Dqt9wYPxFRCmhAaDMs7eOGIrlrxqbHO5KbPCLgJeTXpTG1GlgD5
k21tsVEDPnbgjOna9M333V4eeanWdSYVtQPWj5bB76axZLuJf/PGalAUsjHLisllY2WcNBqq8FxP
sv2SL7K+XqncxXU3qWSZuxlLcMyQQ2gh3xAag1yORbv++yUBzV9GhAQDOUo9A85eyUSEfUVb7Zzs
A6j8kM3G8QcrlU6yCMI3DF+6mEmb6l8xRUY+TfkeoBy3Jd7b6MhMHA8i5vMMds5kapV3yi47xtUL
GibuwNadtUVd3i2kQN4eV+CKrv1bZBXNRxP7H14hDAgnyUp5QZ0JjmpdsYroHvbBT13OYwRMcLfI
Dfo+F528gzA2YufxPkxwAFpfxv7vyfGLuaR/ocN1ojro1CU6xntj0rUR24gN1PMYAfo5+54wXZ3P
aAWWhbBaPj2seW2aAFxmPvwLoGr1nSlfH40Q6kP7jB/+v5KwS71bI7rKUODN9+AU7PRAgshr/jUu
Gk8fsoX/2alCdKrvkjL2V1Q2EBgJzB6pKIrGrzXfR3CIfIcHxkm8eCN9LyrGAFbWsAquSzMEWByG
cHf1txlIZLW0zjji2LWPvuhFQfeIbcC0+8KSHFluyZ0r1CJsfLIEaQegIT6n9qqM8ZziF0qpSIJ8
eBRW+ZqD7IoVU5gJQElt0Ce/3P6KfhGPpgePfypejNGVk7NNn3LPyif7mEKRdwglr9NedytVkq8r
wQMlG2XH2IpGZu2tsOT9Av5nteAzEhMzktIbXLXhx0FU+s4htLjCDffh0w6B2RwiCxtGhQsmQlLq
1lnKyLz9iF0iIOpePuYTLfXuw0fR7oppTsb8yYfjUNPGjMYjNovo4HLDXweNUnwbqtCBEcSxwuji
keLO3jaUTde30nwu2PEgBrJS/XM/ytJyB2262/AfXrxjjN4yrqyFS+l63IGp1v/GLXbMZZFmVVpA
gmbOQCEYLs4Ubldoew3HrTCVE6Tqvq20vfKEdCctNq8gcQnyOIfeSdE3eJ8jyVxxYHaePCqCbscK
W+7RaR4Wgtt1b69hWtTJEE0hh+APsFo0VN9dC22ujUIUh9TrpgyguC0UKssqhed/w6v+y+LzZvlB
/kGuXRX+KK9T9H5kNhzA0fPJOXPA6VOqf2toRYKD4yGDN9gNqT76fbwy8+eRyWZMbYZEsUeY4Iug
5QCb5a9d4NYPBx/A5hs4xDO7w5mqKjoVJA4j4yxZoO0pIs9xn/VJirAYU2ul97mhEQxOzCNsAEII
WCZTgjdPTubgKSVPk4lFowfOdPB+6WOmMLbZX+O5UByVxqk9tbWN70YWTQvysxYBfXOBG/IyDhDc
PEdcOj9fmKBZfRQ7/WjlXfoK+m2x5A3GX1EeQ92RcXL3nO1diOsbsB8tbYWCt0CiYG9ZHOQ7IpRE
etlw1WMiPTlhIPnmckpohMY99AsXMLQbwCx3Zi/ruSgPAyfPNrkYmtJTEgRTg5FKqMiNcGGzIh1E
luXX2fOl1aS9cGyBmUDv2cdS1+OOnobdStdvSNPA/+4jvqWyXTsJWitwhC/xRY7EWLQly3veFYX7
V2ciPpOdMOmiKTpjoGKaAjna95MBcX9GFu9P9/WZYW2ClwBBlE8ec70s5/JslApXSSZLD2AXuQx9
ktptusucrNhQ/dPz1B6s+9rOp1LRQw2Zz9pSOo9P9SkFQIRyll7nqc/XE8W9eGrnxACZ4uFPWxUO
wBaevd+1Hl3y4EE/noXIyCzeqZ4Wu0K3ukAmVoWTUA7V9bLI7+CPk5vTxTpwwbjE15Ry5INC9kFd
44RiTwdHhwV2Hvhq7vDG0DXbiNNkq50HOSMtdN+X6+2FEDax4AHZ7RI52zVWtVN1r6xI5knnRDvQ
xCtZXBWbjnOUDC4PwcNO8CYkETXlJSAEyOLhN7yFr/SKDDpTMAvagzhUIDXVUcayMjyBTTLTo91I
2iu2+mfXjJWzTerrFds1Y3FzivxRadalcRqZ4Lb5RISUfcpPYqWaT6rN0J69ujXEdIM+Y2fxJGWY
eZ6ZcvghZiO9pODVhURs08XwAtztmGNfdjpkoKy9WywWY6Es7EIEuCgSlaYGOyW6o/xMqGdVDf3e
Fh0AJkUPLgmIqadxPp1Zhl5IDxqgg8vARXpDoXdlp9t3tAfja9jD8e9A81lqKo7aIhLD9CDy1pX1
RN/oV0phvWFclGQQM4rrATJYBrCyG2T2ajr+GPY5MCjjUbK3nEULJYz3MSurLywfpC6uthWxFxJL
gUSuKXvKY86M7vmU826ID1kcgJao6vgX/d8zIRL77aWc3RceUDMRqCL698sUPhr9A7ck71DsQBY6
wmEgrhNu1gidfULeULVZ6ehR/nKlOarTu3oYYxtvISE/krQiPGVytlGLhNdjr7emZkiKX7A3ytl3
nz5cOvRc4pixsM2+d8n9oyUVNFVqQTTP1Kpv1Zlkzozj2Szcp9DpAgNspBq7roXRMGApsIJcOa3R
NnHdNEJhuirHn4vUw+YfNN9t6AiscmGN6wsyWuyH3xz3iikxOS/rRVimi90j9FQRCF3fNP19DydJ
NuCbALWxSJEWrJgK2Aak4eBJQFx1x+EpST8j4l/w/xgwJ2kMbyFNZi/Xcdceo3qRuqGuRthnjnf4
QMi6erqRxLXNzfymM/ZFy8TrQwRA+br601aLJO8brqsow1ysI5ZFGYDFPq92uX2axQfOIZW5RBDN
G5QMWyNVJAVOXv1LSrJBVHw2SnbQQwsUXhTd7/YSv+vdD7ojnPOFOcPt7p7HlDl7PV0s8rryi/37
ulPyUVXe4nZLAI/MBTZVT1Ayl49k2fz4s6cClpoCJP4fb+tejISiZTt4w6g0rJ2vHVCKjchDU2op
BgL9K3IWdFc5JNDm+z/XtEhyLN0P3tIYLwig8+FpiGZveY9tvS7LKkcxoCEBFjfa63moXSY+kdU3
K7ww/tqyU1IxN9lFNObb7IPrkTyIbVKXEY2NHyCkr3kLfEuIibDrCHzJEBVJZAbJxWE15Dz+lJ0G
ja/iFfsonU6yPWYAiJZbOea9so31P7G5vqLZbGoR7JEuEpyN6qTOR4lv/Rhj1YxPH1pbzqrmJq/7
cBcpLt0X+778UvmlfBlDVQAy1VN4NAiIN1wIiyEIGAquY/hOTqScj1ytAX913IbPfNH5drUjwLpg
tc/5zl0+tmhTKpaBOk3pXjLC4Nrf/W/u/dWaA3qSYtV6EU8zSu13gplDGc414ZOTTkgmu3WiYuZR
NIx+zsimzOoSoo0xtaWE217JKyizWF+nyhKAt1ivG14Ku8wEvixduoRBPnFcY3hqPt63UUbTaRZI
U/TrR7R8/WWGyNhTIF1y6YbDbfx09OSHl8ChNEs0dOQCeHKSAlXmPS1OQG8bcc7pxI+0u8auQwPI
PJLjXzWEOHhNsFmabzVxWF1PCzKcw07BuY7VWaDM68GrmbKQa4vL2j8iCgGsaMv44aXkjmtlIY5F
rRbszzIPq7DP01dDl3grR0O06jSgeurAZtXAXBfO4u+rYgiyCI/eJfJ6G9MIs4rgsRPk5XWez1/M
knOkbu+Ep/S1iNbCIA/QJ5ABEQoG9pSiBj7nPNN9pKHakyU5iY0J2g560ejmIYt75FhFMBeJZnSh
tqgNDkGgwuhEifDyRPBcDfB4xK9F3Ib6AhibCqA4fb4TgSt0dl2NLlcndabg1ua8TRReHzjDL7U0
sp3KfbXZUXIV9EHS44CtaOfrqjQWIqsJL+WYmZj/mysZJcu2W7/Z/C+gb4EcfU2ajWxFEaLV1nKj
ISwDb2or7n2CbHQObRGTGCCstKUSi0yIbMqlByVMN+dICVl43S9IZGfMsp4blmIg+bWHtl8hDkf8
jnB1NuH84ZTV9xQ3br78/YTnhH3n2Ye+BX6LJwk9aLyOYJaSNdyFWvNSIC9M5EuC3JzSfMelAzQS
iKX5esprl8l4tHNyXPJEMXEHG5wcfs+vVYvsHKufPVqj8MFHOw4xBH9juRTe4BLWhK+BEwV5SGQe
3ntpHKvfymBFZYHFBoOoQCYWO4HLfZjIYjDQJzn62na2CN1scHxuPtBTiSy0r5Z9SA798jCwtDOl
ukK0vk0JoMe6aagjK/fR228GyPTPxyEL2R30rsixpEiKF0jVrRoECrUseTn+awYtFGX77hhZPdo0
zhO9nEV6jNchOthSxAxMh/4WSoWkP9XRPrPgeuHD+XUxgXsOdE5dm3qVlBMZ/Uh/m62MRKI1M6QL
ge5FbbpVvkJOJF5KGLpXP2YuYlcOFRsYfiQlCX/re0sPlfstCpHN37TYrKIujp+v1+EEPAnQb9B6
16Z22cJvSrsdwqHJYOBVMnjW2GRIksqCHdORscZBRPg4/hz/nQWIp92IlUUHVSZK4GI1e5bLSDGc
v/ZVj3qFSvQMdn42HRyLoABoOWMv2+COaCE1IntYy/AlovCC+eR6JQhkh6Phxh5r+h9Pako5Lpeq
vMeHvkyBm5AfgyzGmpp/D7JOY9g4aGubsRFL0jm08dNHau2NrzWHxLQyorK71aVO1CZdxaaPyt/1
pS37e9J/HYHMJ0oA/hXBUPrBDM2/Dt88AbZW4llBaqbKaZvixvwadzikbmo/WI/wYC/od0gMVKgq
fAluCqG5rC100ghMaVLfKENxLJxxiJeriEEz9+zUYHsovzEITivwhjhhFe+vPngaMQRpTKF9EtCj
r5/QULsn3XzNLm4Kmm1CoFpCFQyov7SPxudjrHjvf4LY19H8+gpcetJHWw7Oz2D2CQp2aRoV1qs+
z9QjZJhOKcR3IyUa5ewjj1vyH3PAAy3Rux3TIqUjQiFFuoYCXtsrQBdNuYldtb4F+u16UHBTMi8j
p/wcMbLMgopgT2aHiHx7EovoxVqKVGBDVqgmu5XRJ545vQwuIVEVd2c+yTHhyiGKML2zKbgL2CTZ
e6KK/2al7OSszejqdZxKa+wyJE+ijv7Cu47BJVGr7Y6v+8H4krfVPpEa7+NQn/SNhEElllgpN3cQ
Hs9/f0hN7E9JIb6rli3gwL+FlOlgbFm6LCIHfvBI/I3AxxajjyS/oEfnbrbzF8eU+VL1WrZARpHT
ZoQy6f+xniWqJHQqRRzTTT75Z9wI710sKWs2gGsLZ24OrE9aAopqjGRXfjInof8R13yUQTwjmL0a
VzPyQMKkddyW8P2OWHEsF+c1aI5ZIp1iUhxZOvmy2iTB6EemusX9tR163qqudEkD8q5xTztsSck+
QQkm5AmxYiPYZjqT57qIvIBW8CCmKOKs6XI6cl4FRpZpSjkP/umoUMf7fm0+fSIeFpFRFqlktC0E
WCJv/ibqPAcsP8RLbkXqMqwp/OrhXntgyszORhkvpgqr4f3bJnhe3PSQKPUtxV11No8Hh3Mv7i/O
YH3xbxoW5Zg+QdV+LGQb88V0MsJwbORvPcHUT/npWms9U8xi3TZV3noEnNre/nzbp1kG90UP0/8A
18oqI1i+b/bNQaq++VH71HSkqUYYK8znJYjD35/dJDUT7xXxy+m33meQYVBlI4bzC12Dkk0kEUbW
ybTB6eLzCkDsTXoXzUTF3ZO7lYcg74KcOsi+R2gMnTldRu+vw2cFNHzbwDtFAsIKWdYXYctbElmi
FBlUSWsVcLH/zPQ6ZlFbRzNBeQPHFXP1s1FWYkqeWDBdvMJgwTbOqD9tbLDVoUCBUyR51yvrx5K6
GiDUDWhk9YCbPB2nYAKiZcLV/qYJcIUgno3YZLHgLZdoJOP5XuC5NePxlf77dRzgC0Hd+GLpx76c
4wpJNOmvVOGrEe+C7765CYMBShzdiJPx1ecaDcX6JTq1A5aP77y+QjCzKsNXggxmR9ML9PwwK9y4
Rt63lkJfCF69Z3HBfCHSXUkvjxwDqYbfzZBY2wgGCO4fQC7AkKy6f+jP/ZYf7tglmZ9Ss+cG3wbe
tkU4ebR1TOC0Q3OVOkGC2fuvqoyO2leHQFo5Si4UmRF1qdzVg+Ph84ZxVBW+LaoPuOZj9rKKn9Vr
lpkCnejbLaJYDZcqaFq+cqdRlzytR4eDdXWrd5jlEkf6rD2szfKo3vIaxdzPq7EUbjtwM+4JDa1w
jb03jEdJrt1+mq2+UAjYZsfmPvS/xA70zgky5FM1yDeCeWYNjixFYwZl+P9aI3cCattalSU82bvU
nfeR//dANHAhXZ0bS4vFVrGUwr5eJlw2KgvYTbst5SfXuZToj5JZqpb9jikzdTgjGuPg4sXS5bfH
VJVOUpwjlm0lIIUn+A5+J36YdMp1YUzcMuVQzyUwjgdc8aY5PGuzp+dvohrsOsOli+gY5H4YNO2x
gJjiP0F2LLV8dFmL4CT+L+k775abp3MCkuJ1BcGbw2bgIZThO+kx/pAghRGGAchz2/8vThxwAWdG
1BJdu9brIkK1RSdUq78FJJCNfcznpL/fdeVu04F49zigmHyAOCuPcuR1uvZ1+TR3EBveMPNwtHDM
MStXgiYpPUwVcLiwyM1Z70NBqFaPilAsUXrUguDHgqnn2LLB14JEkSKxtE+3AwlI8v/zDaRp0Ubq
KpIsEHkT0Cd452Mai9DlPNS9Qx15PzjjTLdJoMYiApGCzPUAhbbmWcFoRzRqWOcbkGbHck+DD9hY
uFB0CcKgwfcJzZCUrD6TJyRjL/SIWI3QRL18d1O9RZpAb+9jCHGnM0paMmczJlNIWbwGe7VgD8pW
lCNvRPVYqgAzR7CZNVddeU62yro7YF7ue+j7BEwcDiJ6Qw+EtikRDeVJ9u1/22EwQhu2mN7Nkwpb
VWjhgxVYQ77DnXLxTxiYuT2QU6+zFbwX0Mz/Req7z3FonPJFBoHYgwuhxrsm+MRlU/Gw9YEu84Pk
+Dtk/U6Uq1L5fPyZakM5JHgbVZNdG/rJwHXcOlawdq7MMXhATH+pVtKhphgfTsPdI9FH+JzsLndI
+y42axeY7fg/BDxv3LkuJ3ZIhWrhOYuLuRDnW6q4AOHnAb9uT1ys22oAZBZI4tqPgdpMuhyqiqdO
mu3y9qohPb1uhkcPu42sTuV0HkNri5jx9fgHwRw9bJQhd4Vlkz9zxJ0qFmGdZdRd8wWlXCL029i3
oAcKcoPX10iqv0Yc382w9ofFscjvxZujlwLzDjZCCOkD5p7azWbOi7VCHdeolAKksJv2Wtj1QDKl
ai6oM8RdpfddLhtmupr+SbB5sJT1Db/xOhadm/8Dm553fGdKPycW8aiXOwuFgf5QlX3bxYulr3wE
UTukCK90PF1fhEYAAYs9fR0LQfO9h/WsMLDHVstfmk7NfFQSNAffimUnxdX2P44X93uH+TShaT/v
np6mYZAkDAsTl04l23oEvyXGLxGF+Dl6rgzdjq2hkR5i+8wZPt3VljTwupaNw4hZx1SOZxkRAfcR
6M1NsQyrly9pZdzOJx6sRqBcq6R32Er9jetFFZkrX3chnZbNs5sspsJhYLWt0SpD54+Llenqd+8b
+12do6h7IB5r5v9YTMftxMjdMVJEQoYr6REbiUgF710ROorlni7fJNmuFMVqNpYr2cSricBZWyu8
TiFQo5wP5hxt78B1JKlMYFlfHOv5MtiC+b+9Pa6PNxPuL0OOB/BK4nMF23kniU/Z/EYoIgzBRt+6
vnp0mZDQTnKMSgMThmn2FUjkK9DMFPkX8NttONn+z2HD3GYXKugRwLu/l6ecOJ8zpRaf9Mszz8Lw
pZFqJgepMTxIxsLKxBjpELl0x8xCpj4ZO8sGV0PP4acNlKyJLdcDt4+Flh4qikkBGWg2asyUjOK8
bFcGY0nJq/DSOaNFa8pc3jEE1Ms8Cy3d7HI/sZaFHARAVTJhGfd9UZwu7V5pjxIm5QMNnYgA/dRx
txYVWXDT8RqjzMAJs9swBaSDu7qyaCSHVTfmt8WYr1vMIf8XNS8G6ilfgw8jWZPh03dnCcvX+lU9
WCg6ylUBKr8x6ypy0HhRF62pAVw9TJ4Nxte+gmD4m4UtdvlQrCcUhZlSoWUz1CD4hoU7WF8kTqtf
GkpQAri8pS+pP6AZm4XiK/J02OFlUF7c6A6YG50BHuXMgrws89Pm41BmzJYzH+B20jutsUNg7Ww4
z3xuId5e5ot+ifogLTtQK/df1eAEP5NVFOeplu3IIOIdU7r3mGJ7Ciw+W33f4xBssMO5cMPL06hM
xEnjFZBQWx4HHTBkUOBy3N+g+Poeyle53duuE0hkofBNKObIqlpM6KBOTTEdbLKFWnjSLG2if190
oKxGhMxA1eRmlqq9nzMzmRiVIU4yLHN78bP1n7q0r2JUqhijwA8m02+jZN3+Pm9mEIfPWWAQPr+q
hqivexI+KWWHJsgcYUK/AWLhwG6nmjC9AZIokuDarYLJRXaTnZasQOFD5bkCnGGRyGxkEm4z0UEc
6wtwivPkMQrp6E/+hFQpkyzJuUql1GJ/vlEeid0+5utup3WjuwWo/Hur2tCoX7YBkCD3pVPkh6b/
T4f6A2byPyDKQnPX9q8Se/MsMwg/U9b9qizUt8ihNaNslzM7WZo6/LKn0jGi4M3BqVCm+lMH4q+r
+8okSPQOFB9jMy6erlZyagpYdzhvtefXr8nqYxOrkiIcINcVg2fTdKetKnduAlTG3zmujT8t/v2d
G+ax2iZDV8AnXR00gIcev9b6JTIfAqC6wCn0IWXm9HVgtLNf23ZuRwgopT8BmCI1uKsgIWe56xDF
Td83YzdjQ/xCJdKQmGj/3rDGadBPd9UxQLjj5DgIxnLnkAHYAX5GtSD9fGVGCLxnzV6eOJRdr8vA
z/2vlp10Ymr2BIp64NnpvYkwCbCGnL+hDeoR6NzX2kNnP2Gb9wshNtai9kLlU2NLMvsSe7EiTU/g
Q40B2fdr5YFDwBHFsEM4fpeeMCMc97FkiB7tPCW6cmXQGMDkxqDEM864pQ78FJB6xRs1YnR3pW5p
lspHnDTurmrj6YIwOVYcgqLtOia+/yIki1AfnXrdzQpeq6p2ckxQ/Y/bYP+M/Z7AzQjsnAbYGMEo
ycD8VcSe94120onJH1p8aHD4TAcdVNtaGRDoIknORY4/GaHlOqsIgWVv7FofJbuGiCPItioB/wO2
VCM5VDSG1/VrtXM9YSWUwiZS/qcP4UjobDejMR9JTdrr3T9ZVoHCB78fqklmBIidpHsjzjy73rdh
zs07HHz+MvpqQYYsn9c4rpZX7TNa0grspuIW2EaKLE+nGPPmJZ4wwQQFAuGzTdAKDqeqmzhaV5O8
UAlN+APZFCF4LslOPWyyXqAFjHdLnq2U/AVscDIbemErMBqUbrocD7Kz5MX5Md5NJ55zbw5tGvQ0
O7BbPDrexFAOZ0lv9EVkaXYw1mWLq4awZt/BAe9QcxZRjxvalUR57YWVm7vbASoBL0t0mv0fHsBq
JIzBMkiuyVysUz5g7LoWoyAV3AkOdhRb1OkGOEx6+GPCFVB1O1Fi7c2r3U/cYHEAnOU6XXpOGKX4
FxX0mxvEB84OQaFePY4c3dSBMHXdXrrmeqVmIggjJbu/OkrOsDTNlwlHiGoRjGYAftpwffOBCczz
h3zMGirDdpiwMDVq09L7YQCDX4mOb8v74aNLxFqbPYAu6orsqP+wmLHNECt4gYbKgWxZiNOxb1My
Sux7ad23YZ0AQylDQan0ORj8sAOYHa598rl9lLRBqwTbyaz1681vho8e2PtFv20CY9qifXctZwOd
dY4OFRKyx+zdtPL5ICDLUpIpMq5nwm9LWY/I61DxNRpK3H7VO13MCgNllyh2dvMrrTN/U0HUOnjt
EXG+mE5WGxvQIHcGDfZ2O+nPwf1+DdLvfPRNNhdFrt9XugL5XgTBLbwu+U18xvciLWvCfKfwl/dL
FldaLugyfrd1zNvKq5thjURu7ZMOkNrPpVM5QwzhpSh7v7Y2VSIQ7LFbRx3WARr7z651spXVC42F
1l6PohNoe4gst2YKuJn3ICqYvQhFIIQPHRdO/bNulUJJOWjm0Qj24qsQ0INd2/tWeTJAIOP/OEhT
UCkK0ZJHsWmFjJNoGWXzM8eoRIGxo+Vewh75uR2fCRRpk/QhEw2JmF/Fhs98c1Cx60HsM/kyIOER
IUiZof+vqKLVkXdRZM0GGPEHT47rGM5JLGo+VVYCnNjH1XZEV10utCMU7OTEXUWxWWphYUOV3Ub9
IFt2r9zFakTay+b3JIwisV5J+BGfg/v6EsE3l6aLSxSBU8WekDRvgyAyCfus3fcEBXEPoKyxq466
FHOb0o31wRyf+YGWwsg0pvCv5PK8SCIL2azBVBp4mK+tdWe3lyCf8WuzMnHbiv/9ubNtRIdXrPkt
w5Rc7+GowtQgZrNVyzjfV+epE7vNX5rMmnhugJMtRskpoQIDMjZ+JzYVkfIc8Sbka7JHobSsUFex
7zs1sZRvrFmrxFuCzWtE2Eaxm6cHvaevvcdXDhEspaVYQ57jqQQfUYRV4SnErESi9RoJC7d0cI5L
+2iXfxsbS5FqUmpTi1MaP57BQgTSPYwmc77nU38ZLjbickHoVd4ZKhn5xAiDFaJTnVvZHuCDJTIF
Bl0p3G1/BEHo8vop5ZJrN2oxrVtD9EKfiTHtXwq+VDIFHLZj1yvxYV/rezpv67cYzja0vzyf7WmL
Rqw7iXEPetKGvkyyosFQzfBC7aGRYHy/ebLRIJVtvNAZCIzIjbNIBXFtyVUjZGRrWKQG5URVn9OY
wXqiHDHCaeuwyWPGNc2zz+svD9tzSrpfjX8unKTYkjAmEwfxGu4uyJ5OOn3yAqjyAotWp1OFGOES
M3faaRQh9E5nDHG+R7g0/ADv8eEpfS9RHkW2wndPzcVNeLgV12797UpyOPnl4Ze98lASu+PXGUGG
kBkPpqSCUd6vpw0svRn0jirrw/Jb/aOjbmXxzOviMNQZ8EtKGOR5dVvU3y6sLZyfeEj724sWGtOa
DPrRPLLARiI89FGBOV8lJohz3RVU0mUraj9OTumJc7PeJs7LrVc3ZZafQAsGFAgoeM8wdSdR9tfq
8daeJOfIJVLH/3hjuBofbD76CxTZuL+lOpIWV0LFelEX4KtSQPyb0R6Q5erHGkhwuQCXq6NaGFrI
xA5rzVoEYtpWNOL+jwdHKM332HDbm9rF4Lk4mnDseaXqtSFHEPlppm4cGYnWulmgsb12UIv91qtA
Sh1/B6dBFhGcVb2Z5pl3Vxk9Ogt4OdDE96IhMVXD8fi/fX2xruB8UP4owKkgO/jeTxj2AuyVm6GU
8rjMaKhZWcNw3UwHUDVnYXseOsNhvEwIJqivhUq2/D+bXTHOHCf13VcB2qKu3R2NNMckULby+AwL
jTd1NA8Mm4LkkjKc7xDGVa/Gi7StF4nYdcihvrCz6fqYiufqBWdmq9oXQ9za1ZnLKUiiGsy4rlrX
89Kl97mHMk8LgBLvn++bNRMlXquYxbQrZw2ecGcjY/z2kwhhtc50Rl8hXhXhjTIHoofsLUuO5mEQ
L4cJICV3Xl3Zp3t8MgsrgCIDBG4N7srT4z9ecjTYRj9lg7kEu7iuv54SNxPE1I0HxKVpE7CbdMb9
M5cTnsNWlOY55YZZhzEkEfZd890YrQmuwuzfl6NPXxv0Es1UDZUkSuLm93y26XUWC3KtSEQ4Vr6q
lIIvpQBVpMxqNXfDv+2KiDL9ZKWhcKk8N36hgTbPA4t0rYhlsm6Co0XxulmOaErQVjxgGp/2p6I2
4jrsfxVwWVKd9Yzj46d8UDhqI/aEoHli17jOI22whWtA79VoVlsglsBvECejhyvW6Y+/LOv+DQBN
jSHtomsxPkcYk4TmzZVAjAzDxGqyHSxW9F5SK8rzjKSQD687HT4nCy9GgbNiyuWvhqF52HbJ4NPY
D+tdoAPJZR/SurL1s2BYkCAdIM5iGS28tc2UloNIOsuf026CndMuI/GZYiITGHCgEgc4+27QhIMs
ZUp5UOX7pBCD8+dfnhKX9gONvhZWO/4t/izxzgeCKpqODJRIQ8Uv1deJFEki/xsFLnUL1UgbUyAA
dT4Id3/gsUPw9s5yHQm04Ck5eAdRnHDnK7d1+v3qINtGEAXPdYFUH5XUk4uYChJyN06MSC0Ed9Ej
UZjR05kV74QTvEuUdXy7I+2GWa/2rLUqTnuK1aAdHDG+rg0uNAcMcT7eeW++IBHpRsB6Ba3BXINF
n1aDODYNVh1OmfSVsEGcVgpph9dPAjBoohRF0spJ0xo5b4amhXDoyr5zDMn2GdXyV3BDKatj2UnS
qW2GW7QwkDXa2AkTXW2an+7S7qdDwsMHM5jhMFFMHq8+u83BqJybvflwoga5qFbmW5Rh74Vd+2Br
qyZjJWQAvm7QZPLStGrIq2l5IvkW8nBm41Wzo/TcJ9ili9GbC7oxhWoZATHSSuq5skwjBAskSyfq
R8ldfEK2wlOrG+jA5FeHzaLlqsd8dNyZPpvq6qcNqqXk71N6/7B0oLXFH7Bc7LHFUnFKchZd2bmq
bzttoGRNM1XeFojWwUJdn0Os4Yh4LDVr2ee/KgLUCb3cPe9uQB3hscjeYbSyeOO4xTaQyXY08ODW
EZC0QAI9bmoDXSlp3mlGAGODekBcfQtGaQuC/4OvTV+JG1w7x2t0L/FaCLL0r8oSrYjsaOgkgmJ1
MnFG+FCveAftzi9I+zYXVayngAW2xOpgbbwmKIr0Innfta+FciAaUlsaSz5AdnzugWnBf+yZmnWJ
fkM0tXhzrcWkZKIMimwMCg9nxig7utW9i6xHiX8KZtxRaIcZmKaZbsFVVnQJH5c60yiPLvWnx0p5
9XaWjv86FvEvA+ShYr6qH4S57brmB5wXeEXp4LEi7LmgX9wEuBH2zwWWplY+Q64KZcBp4GuUARTQ
qpnJRcD8TsXbNRF/IkeqjsN3TKj4D0ibsK4YbjF9mNCqcbPBEUCXrJtnLLQSafJns4iH3bNiPOtN
lYACoD0oJhnvuYgZbil9/tY66e6OiAWYGGPHf21yWThTD6JZkJ5mYz9q1tC9PpaqcoCuFVfdM+g+
ws39jwkotp36XrS9Mi8hSfT/Q5lfOgaiZreKxrjK++xJz4nz/kuOUqKciiEH4sCVQo+H4zncdFOU
aXOOtD1Hz7XlwSbFLmitjZ9gOYBiKHWkfiy4kL8OBah8/7MZjvlW2GIHWteXR03vshQ490V7BIf0
0ttt+lMtu42ObUeBdcRsefzHM6B254KKI1Q5TcSHCpblPoLFMAL1r/UZ9bg/tKIi5zggwnp5dhY+
FSrk8uB5emns1WuThmO5CdQWD1v64yVhTc5aTnZlPJH7asIbrIpmtQV4/5fxX/8WJ6TTSeHRqTRW
JHEa6lhgb5De3op73KBDpjzreYncAwvh3g4J+qYmQeel88zSoxZipyp+rdRrFZGCxX29/8mQDfQh
ZYOsAQ3H6Rl8hHX7tZHPgEQ83lMqGUPYcYO4dt7Iv0h6wwbqyhPaPzjxrV5f7R8+kUeYiAJ4rDOV
1GgNquad+jlqXgrvRkkwEeS6ztuX3r7f9WahQXcVGGmiqpvOoHyhJMciK6y/eWqThvXtKzEbPR51
VsYSV0LY/iPsulX2Zkkr3TxUmGzmkvD0IgAq3J0SX0nENaKubjzuGdegM3EjzE9wnPr/dlZw55Gx
YyAkDhmIe3Xl0kilrlAhaZ7PdK7WvmmVnXRZdZy+1JKDxIqH/ezGbEaZd5eqyovPj4zCQ4PvwBUn
Pd9gS0fi+M62NjW3PVF+462xaTxsEla986vKjSfuy/AQIueVy5ehd2AQrkNerSv35vPWhai6xgDH
mWxPU6qThHppQATA4N606VpoR5hz7C03JK5Q25CLCePdMZCmGuU2/HDe/YDQcakx/yNzh8HrfK6t
TH10qkgEEtjiC/3WAPqO6gFd3htHVp7w7JqpK0KxfIP5qPZP6GMLiTMGzMNhyVi8f4mg6VIJA2Z7
GyL4j/NeCPDG38/Bu/RFK5ZSt7Lbvf0mNYZi01MbIgNHjtBNptt+M/DNA++pH/6aItbOo1p+eiTA
KTJl6LyFmbGija6l4NXuxK9K0H03KfShXfdqOlqXCOZAZn+ATkSynE08GOXGAorOnb/iG4bSqo3t
TLVZhy9fr0kixhDzFT/RJSoaY4kV0Bv1sVvGFpPWhTI4Z8T88x6NymruOnYQjsMe+lhLOG1MgKtC
6lUm9DAOdD0/3xufdNsRoElkHIWuRgI5l25KfWdD59Q07cIKmUcf07bksNAsac7WwK7Voc5JR/xS
0q1hwX2Ot5ClW1iZLqE7UVPn9cS7QYXLwUOZkcKi3Qb0UJpT4Wxe74/nsw35xiqLQJva5pprKw2r
pX57lNKN0RRjI1Nhw+NczDry8ELxOpmqtyGsFdSzip7ZGbCDMwQi2z2gPAEJzpitC70VvDbNS96n
V6ZqOlqBSdCNqbjsdLwL3ZLcVCff/WbfFBQ0W1jQuGlRlPDxfvJitXGUI3rpzHakcF/3iqus5fSy
Qo1S1FdUe/+9XJA1Q76DfQWsLSoUFoa530fu7ZVOjeGT8DW04fpkcf4N2HVZks02GUQhj6EUxkq2
30z8qXVQhwRue8TsyO94mPOBnSXjd+GxITS/N5908/djeA0sJA4CVMH6EugMnwaRLU0y3f323NZP
1Wl/yD5476w4jdbCSgXdJpgfBICOoUtZJp+sRN7cOj6dV5626/4k/Llbgkp6YqwvaLv/Puh2l/lf
6N7yXdwg7YkACQ6Ii5msTYqGVeWEQLrE7JRRMO/MnAfrgYbl9E+eStojf+RSyXi0mB23YTDFfpp0
nTZ7wJIMiFDjla7pUbpAkTWUBq4Slz430ANjIHGWUd2UOgMpge1ShZZVPA16bF2KZhpuSDIUhvlK
OoI+qz1BqQb5qIYbkrjVJzD5EgvBmqozUf1N3NabJUrb88qVnje4JQG9S51ShKpDLZOGJ/5tbhQN
HKUMbcJiHMFIyGOXTHQKoo/KIs5ciH0F65Fv6LSgGkZIhJgsNLrXYq2CQAMOSYpj4wtHStc+McOk
YsHsSeIIurYeUN7h6Tg1PS4rhtPlITo6PcHYN+6KJFCkrhLJbbwJez2iiyPVD7iSTdtV4/CWq2KA
b1KFYSK7trACJYYnR34Qtm4KPHaFDINL/DM4mPB2aQ0OpOH04PJL8swdXRG4rpHWpJ4Ot4ku0Kyl
5kegmukSbzTnKhiNv+ePtFO7k5jxqCI9mjlCAKlhzd/Lgbpi3AFvkzJHoss3dEdlsYeu5xr4Y4Ca
w42Xu5BgMpyg7wYuXH/CzBdKSSQxy5SHL+qR/pbhBJBIHzVOyjbJUVImNZSNWsJIopqg/AGwsJNL
VgcQbHQFrfLx28OjL8M4ekB60BtVaMYH3F5QbrPFpDLWCLxMUhQobaeunjmOcMHanf6dNcwuvUTg
0vUka7FlgEoQNNoHY4CoD/Cd+qBsKr2wxDdi/nHpy+tvAKGtk/77baNNLEpelQmlCx11mKi4NQ1g
UEXiHQiJ/hSMG8TR40we336tBxZHbKZY/Mz7wN17t6YncESoYcvaRpLkQvpwWwZBgMRMwrYxX1/n
cfF0lndtlqhGT6LGGMeJda6Yknd1H+Ro4Bb73ZM+QRE8zGNIs70u/0AjgA3ir4T1jRdCZV9FD6Z4
cpCPgw7EhMBdqeJifYiNieO3kzBhWaDE8Vwk8lzFMH4sds529VtIRCMg9bwlYefM3vOX7/gJegXd
fEgWggzA+uc71/3BnTtHclf1QpfWcyyGWDNZJIbpj8pJWVt0Nxy4BgoZ8U7fknVVTyROO+rdHnx/
7NP/JMA8MMwC+j+5KSaZK5YgA9ykFtUq9mfKg72xNgFT+AVkEZ/94cRa+Kk2llZJcLU9t/90U9Tm
+Irh3Xb2j1ma2nIyLH9Ne2jwJZYGkNbQXTwRseDw+9dYpu7sxYEmQf/3uZYdnOZr8fHvbLRvOt2W
DeK5se+8eFp3/1PsRAn9zeMSC7pkf3TrYx7z2aMSwQFC911RioIRhV6b0f1KmX3BZBG2eRMoi5e1
KblnnxZW8APZqeznLa4xzQUSiuhT1c/TSUDIAPEg7Xl5+oAlVTH+WgFvCBkq+pbqDXPuTKV7vldl
7oXGJj7LFTITI5XA6H2/Czxhx90eHGjBV482N174gCsPgqE4/PBvBXIyabxYtDra5m6WuVN9BGXK
WwgwObB2ql0elym9ix2/mnIinPO79TL109Vs/v9rJMZINgoA/F17/MGh27N9ds5LKt1WMDeuRDe8
cjMsxEgRXJSJ+HRrVw6NiU9KHwfb2/FOyBgTAksXj7SokSF1KQVv3maiFTeW9dFNv95QblPm1aVK
zmUl4XWTRcRBcEh4ZrRgC09P9M/P/Wfkff0zgkeEmhUfBdstYakvnccvkAmWN2n3Wj95qCwKtQYq
fGek0f5QoboUJyU0EEELlLWI2MPHEHX1CL/kyjV8YG8ZKZ4gFnHTBQ5nu8gkh+aRSCCfn+XZrYz2
yY7X44SQIDGEJXD8LEQqGlpX5kiAMDoyFZZ5FmmfH9vkXL/HKv4wvmvdS54+q61JgKr/FcTavMdr
P482oP0E5SyuVkW1z5b4Wj7dm5/ubr2cKbR7ZeFWlCJW1dR0/076DVvyYcUbBR0AxnFZLOWxPKyj
d8+cQtMBN7gHyNdf0sJNoZRRGy9Y4hA4WK2K7caGmNzuh/MwLLeOuHxd6Ihc0JtKpgSfYwukq41N
HZ2u03JbOa1Cx34EmxNC6v8Q7/Q9jxUxeiJvdp1LYMu/F7/aE+bXjVE/CmDf8+bX8EW8xCqW4FJA
uYcCifqRZBuVvsQ5ZpV34d3Tf4lPd8x6W1vy4V1EPu29FX8hOwcsdR5fddD+gBH037Qex/HndCaB
wjUJElHIBotIZx0yKyvxn1cZEylRy4yjVa1VIn8aFhluSnuFad9FQa2LaXziNsxFe3+ySLlQ71pA
CNIBW0/cXxNJoI3FQMByGaIzrlzRXIx2zC55AkVFXyJ1CYy7dDwScVycG21xcNV0YYBCm9IUGeBI
T/2N3Bn5BQovZl8yMUOPzNs2zNuIWYcRS96J3aWWpG+zdjvXo3JQQE4buvMNgDgl5P0zD1PxLGUG
v97nphPSsnfBo5Cixy7fEW/pY4AvbHutAl1/mZRIKuuxD/A2b8dNEjLi29u0432IeTXspJHofqe1
E4BvschViQXOx9OqwiNzen0ozSuDmywdEgcUXv577bbPEp8bc5SV32nI4UzJ6/jOLdUXHrB4Wnnm
Jkjv/OOGCaFQqODE2CHx3JxeKzZ0u73rskm8RPA7+3pWgznJh3MPBv1dBm4W5GCjH2Wwxt6/fI87
iTGa2LuYR95hYPcHiJWo9Yk9tS3r8kfWECOt3uoYMeHyFu7taptd8COaFCdBObinqNy5U+iG+fKN
MNw33U0ZV9CYuocPeCohaQtOpCi2leM/EZU//IX9mncHFzCRMlSALIU+Vx8IelfxE19y2GoW96yy
Dcmmdvmz9xJ3L2NaeZjVlFVtMLgDvnRrIXIioIaouihb/TNUh/1syaqL6Z8SeQek2F0uNhEJPw9e
f+wwLL6JEoBk2EzIdLFBqAIxtP0dIf4qulvdMSO6zubW0yEfUdsZWJs8PGoh0J7uIw2Cb3j6yBlZ
mMoXgEGR2su+EaWBCDniIc4nRZtjZLqx7lIhXQSMUEoTCP5zvHFKB8JdXivMghyQItK5OKS15s4T
6UOBO6Kq36Cw4BFCoieHSoydqDFwWp2XfJdZNGF4BQu7tR9ZFtnWTgpu+h9oHywOq6X7PYSV63Ut
ETH8wreCTAY5hkTjRF5FtdL84b35lhrST9/KkQFzpVh+BSleBhqISoyG7vuGrKasxJ0uyYuAT55l
p4Dg1wdWfYlAo0451XS8fay7eEPwdJa2pJVZMp8akbuQizzZRRgqBGDVS1Cwsb3rir3KCeglRGEs
MLJU6ubD1IcgZIAFtAib/at8YOWuaI6NtzKTzhojL9q9nsXImWep4otUiGD/VsQBN7FjegDXwFnO
+IdoPhQMnb7YdLmt/igdl+Z9qbjNZWoCa/0NATZi9ljfnYjgjVVPcfvIU6Qft2Wgho5+7PF6nE9X
IH3HCPpcwbr7HBUEtYR/kneso2YIUf/KPrvq5NnluqHdMWwlZFvDwLPztuU7mBEniX0mhQ8XZnN2
2LXqzkFTWP70ww0fyJGKv2HHhh+a2gtXIu/M8McuQJwSLwOxHcPGutCH3PKzCg4LtFGqhLmsHpfc
PGBO9OoL8WRHVeEomWHVjR8lOz9b/1KDAheFGpsy3UyBbfDgxCR9bGQ9HP/CAC6x5ZOlA5AaquOw
V0zj8soaFQZVa+qPvQhky/co5mSKOwlJs8P53bpV2rQZMQosQauGf/Py5L+8kMwkPXen1112Ej/N
IjOVulog5yX14a+mPgCUUh9yRDZc1OJLtMwwroIs9nZ7x/FDxPVL1t9L/VSY0vLIDjmlNIWYUmnx
4AY3KmWdAMTxfv+TcuG7BL85u+YaeXuGAfJSRQAN10nN4Ako5zJIVRypRI2HlUULEJqc0/sFgkPM
rdqMZzxQvXT9dEk0n2GTnAb/gHfzdzco3bBcd9EhovI2V99R4L4J6NysPFOug4S16E30db289ofM
+6YFZ92FLnCsFXB6OLngRk/yrgqISOOTNWa15MZhdxqyra9+eB/M/b+gsHQcOz6JkIn87qEx+1Se
GSGYbZJX41QCOul+AvD6tDrlLxsPYuf/lp6Fyv8TNK4TM34AbvliCgZkvcE8gqxwV98BJjAqCL/c
YVbXRBpsgXKCjwv8XSsdwgyK4t9kRwx+eW16tmdz8t68qj8Jixg2N3hByGQDtwEWOTjTlOfvfFzj
IBwbHWjluIVsBiMOFpMQjID7U04SDx1teBngclWthdzY/5zl/mgEPoguDi+1UsYE7krXzXuUasrQ
pj5LtinfdrHExAhOH5KDY3tnthSK2z+9zg8W67TBBRTPAce3Bj3qmOKidsRQlI4oqQ8WEyF2va2j
1lnSpddKGuMDy3mSTQZJ0Wf7nT2i/k6IB9VSGqzwZf1YysKWkk8YaAYd7MuVPlzEcFqnCRr9qntQ
wMFFbEC22wWn3APlxZnS0olcEL34lWaspnwGFT3qA/eIf4Dtegu5sMjBpDLbr2oGR3OwJc56/giI
gOhKOsNxKRXXfCHF9yXoh3gK/c4mgVwdP0z64hvvheGq/vdwr3sqRl0pKfa0iyQAXP6H9dEQtgt+
6rzY3edsWYbYw0KWtu3rKnUdVVAB9Rlj4otK5zHe1irSH2SA4ZpQr3KMb+WjVquvLSJW6XzkKWFc
uMAMKBspzYj8N5y6d4WK1rIYmyq79Ojezr2rHjw+0in8EIWz/FbQuAWciOduTXSnWksL4lfoxd8s
vkuEiBqrYS5Kux7r170eAumwBW1xlk61IwAqOPtmqXz2CDLe9cA1BWfdgj7aGpibYArNpyWR86v1
PysP5bZgWpmRfwIH0MX3uSK7blDKbEKGEqdEhJ7iyWnIWVnTWYMNF5jgshdbYIpRLOx3qE+sbGeu
YKRPcT60IEOUdpUrw290db+v1i+0W3Ht0p+OgpEeeRtwAYVGAjmobtnU4NO1p/QaPdD1E6GVm1ZY
rQ7aeXkUm890M/SIloxvpo1u+mwHTblgRSuK1/9FX53Hor20wKSZhpRL19tUbsmexdrymgB27cSo
F721QioaFmL7RZpu8NT1Gpet0NrtDHkqT9AWfjIqJVv+kWQYvlSWbJwWvUOPbgu9RcKfVoecaZAn
yg+D7mwUncif9TaTpdHMDH+4K9usKhlzaDmbNEf2X//QCaHSTmsYSYyznmYtt0G2XclYuEaPoHKS
PmZhTWpZ+iPx4Djck1WhtR7eg8VWpi08FUCP0zKqS1m/te900ge/O2TC+rc0hyvtFWA1aEu99A3H
eoAjTIXGhO5UX+a8CUctNMRRXP9/m2/PeLCgq/pkPyFl6+n6OcTmOGCM3A+hfQEgazDYiNtD/mbH
6cAnzTZQjapb6+gMz7myarbxavMi5P6WYiQjDkwfKQIbqTrcgWvp+uZEOHyaZtWH7b4mG9ZzQcRG
MPQKPmtJJNxtiXM7hQd1OEH5WPza4k3WW75WqFZc5+gu5w9JahPvD01rrNi/gFpRxD9rWXK6Geqr
gzRA0lOvM5hVUjM/G2guPFS5vyEFKVuEFs7ISWkTqwla/bwEy7Cwop8oN7sUPvuMPzo6FGv67rVJ
gD3faATXtpmqljGSO96bz0boRNEey2aiNBMdS5wfTEmzroaSOkEeJfYlQpKAR80xRhV2SaLQ6tG/
iF3F/8gVsbJV5Bcdj9e/EALH6ktJxjlUgUxdHh0HikcOTuYWnZLxrtpc6233WIZoeZLZNiCTOOH5
O6SR2BWDfEDZzcD3VXEaCCFVfE5JHmGI/CjwIZClqgZlURoFidPxyqGmf8vOn4joz0K0J1IKs8/5
HBu5mx4yEb1d36bGivYo7X4fw0c8Su2GcndYrJRPSfAT5tpWI7sG63NNQKV8bdD7ldpYv3SPZrqJ
7Vtkelur5tN2+WUxauzws4yWu11tfqleNj3v9boyGEBZH6myO2POSxzgWspkUOt8YiszDjW7GBau
7OcoCt9F01jWNvFOD1BUbHt7I9olAk1IOZU0X1q+yyP/GneSZC9e2NZhZafeAOHL7CYJfWbC54Qt
EN9tPvZhOMGQEYZL24edkluuJiDyLMkcYRMPtF91hhM/nQhwHpW2h/ooC13echr6UfraHi16oeXC
fLMx3Z5h/szsxAmOxSXvp52C82ahx+nW4NGjyNjPKG/L6sM+lQcvSZ/EkTLglkZusyXcOH8G+iLh
c6E/wusPb7F/KwDprgE3YpSrY69jgzcvWdhf5QmuVUbulz8xITmSYFFTUCxdTtWeRPhhV7fW9X+4
A2+OefJxkfph2BY8Znmso2jaA1wCScgNlmVD5tqgn6rbgqeb1dHE679aG9yHXA476WRMNGg+Un28
Q6G23rkEl4YYcl1DZuk3lCd62nQiRMgy+zpIonWApKHGw+vFH/8NwKMguZElfQkKhzhsWKFJe5eo
dYJyn3XEX/kLzuZfpPVzustEw1lKYJ0yBENVPJ9WynR4t8aMuYYcYfZ8+Pb1lXnVJ/FNW7ESpvrF
oM3jfUHHzSbRK09t/cHLFWLLgx+zA0ljkjThXUXqdJP11NR02qEVlJkqDxmCeQJ2bCUwB0GoeCSz
hwfEgv9sOmKLbGUCu9fXVto8fVO7plq+GNVZTW0Zb04pUMrs1I6IIdd58J75FpgRqgRbDJKGFsFd
zL7N4PFA+MUXiRKdpH5h+T5taAlMZP/QcTEDVX6VOiBVt+x3rbCimMUxFiD5ibPuXw5RldSJckxr
EQJLP/3UhvaOApGPJJrotylysYX4xOXt84e4Z5iVDlQL9GaP7pnvBfZvT6ifyvv9fLI6tAc7xuIl
F2AuFPZvyW/bZnsU4sO0t3cX24iK1jduoCO5Sd5Yl9uklKHO7hCfsV/oIyrTJ3gSIRrOxhsz3wyW
DMSA0SiwVnQViefA2KXldBCvzFLhZrpAUJ7dNkGgGtF4aCImdvDundNGnW4WiD/oh7j802h1F18F
CQfvMEqa3Djwhz5ZiezzPotArd49ibWJvpOtqhkj4WZgYAM0qEqNlaRKJMYztxabzecw8AACpF7D
eCnavQWAjfS5pivIULMwNCrY+dTjlCXNgxDzpj9xwuVuA8h/NIaFOmSyzNpt20hrKizmNIcNpCxm
On/cYTVka5iTupg6iHy/BJ8M1IrAIYe1sEcdVdte2N+TP9N8TQwq5d1+1d6oiRdFrRUvV59YDMew
QI7C4jUMSx/2g50akf3kzE+C2n+Up/HhMEkzHCyxIPtxLV7W7Dp8a1UWOAhV+UeCM3Py/UsgzFdm
IXY+DNaOUhu5a/DKejXIkwWR75/btuTCq97G72LDaWl2FwgUvzkM+qxCemEIChy+7oYkr/bDozR0
gtQTIX8KYrsV0P4N89Nj5N7ul0vMChrejmXR6l6DS1WoJJ93TCh6BJGTG9ylcqDxTuIq5zriAqa+
s5oi6ezE5vKiiKuGCKMQC+QhBnRLzd7kA9Pd5dABxr9eo2dIX15kkYCchYVvf5Ih7SNI6omHWtqN
LW7dDw5yDZZPeL8z7twt6Ub8Ec7Bu1B+LQzbvqqAOX3YsLkDD1ibu0sgegmapqITrr0FXIEo2uiU
JQt2GgntyDvBELnVIS+WHkyyv7NfV/3Mr2brB7YcKtwosIwIHpmLVh9eYzVxC3eoAmFfaUE1TW7n
gOlxR36DUDbYbC1J/ubQn33k3z7BkdQUEOwtM1nrXj2qage3WKdoxuV0VAzYNMV8tmUuFVGbKowr
29Z4TLP843e6EKGmoCp3/dQBFuUT3lKTd9ZZyRBE5Huz0c6tQxAwyzYeC7/GYRilhEHp/1kcyAn9
+s/a7JyIuupTrRi0KRsrrajnQNuNdKw1ruuUI+lDuwbBx44bbjpFaXF6jMdxbSGyEZ/V/2RI3xA0
+A6g0IZXFzSFnmXqrlOrDphTlek2eXuTCrW+/2meMqDU/uuerIIFr0F0Um7N7pMPFsbvOR8e2ESt
EWnEpYrAixTbHVYLy215LmIn2Az7FQo6hNx5v1w5XjJwWB9XZGREWB/y3iZaCWR5u+cktyx/IXhX
FXhBle3GJ7Suk7tS1AlMtXMfFvEPY/U2F5Kw46+StE2Wu/DJ9cjVza1mM69VU2cqe0UeVkJaqUxI
htPm8Wo5lVRDTOeiY4jB+6SKmsDMs+XEZk3RYG0JShHn+1/pmh9xiFWFsvjGNeICqDCyysPaCbaX
ayl5thp4ZaOmdnPC7bpig3wFjJiKbdMmLoRniWS7juhX2zSoU+XUiJbNCxQYn77RimiGT5ij3hMJ
loKdcOnRrpe9HkWosAlkQR0P9iqLsoN5GM06NfOt+3iVP3zkGuMhQT9+5X/Kq+nw5U/kvZG2eTaO
4JQ0SPC5sVLPgK6DgthVUjon4dtB19S1kNZCa663Ve37zD1XG+zoOBB167JV7Z1WHRFbCo9jZV4U
Vm14S9oaVN5BVrilj9xXgy7kt02KUfzL3YAFPt+t/5BMK8WSgJRjgVmHwbxSRnELuxvIGkcMPKSn
q3u49go+hjvGipEGggXqoZfQ/I/3UuV2e6vRHKPJPWM86ADJEtdIlzx9TPZVwrjjjRAmkdCmfQuI
MO/Ow/pm86cRiqf2d4V4fKSnZcnCBj9fwSqLBQPygTYb5AKcyIlou8KMhO8zXVJSnRP9la4WmAug
Vzfg/uK4RtLX8uJNzywyO3mgMH5zTw0xEfRmU28WmBqDlAhYdx2vmFwhqjDdARplBLax8kD4qRZF
PspJ6G5/GJuiGNmqRCfUjnbP7YqQbnc9dSu795yyQxSJ/kUEtqUlE0H0hC/JqnfwydGbnKaURDXN
0ldKPmX1dsBIDv4W5JG840Fdtit+QAVNaYlQxTXi6LTnqTukczzs2vcUCjnc03wX/ZPtpH1q/rS+
D9Wq+P7eQyrMSvbBLfJKbzgiP5hlkU0hU++joqWdfYlTu/vTSo/e0Fu9hAQnlhvg7qBSg2+fYs/F
mH4GhR4EnyAAWzx+vMYqDtujTdlBSZHVvlhrd7W1hxA2rOqkvGZGx5M8yKVMojfh55GGfstQoINr
/Mp+eCMvvDCVI2CMIvpkVtRsxFXbAclZmNR/7JSNF6nSAcdwqlE9AqThSvtFgjAmySb31Wt/06Pg
/xzoqiZGerA0XpN7IN9vuf+yI0oqiPNSa2S5DIxZiFlf+gMC7iCgfk9D23F5AqyABPJImzULSRhE
6qmdjKi2Z1gxXCeYxIpTZ6OfWhQskIcF0zeO23JA3jE52bfxuV7d94ENuXTtzZtLg9iy17QQxFTa
2tL7fKXcY8FMeekv3SAWy4JtB1kniz9uyzvZXBfyV73l5ciCjTIiX2Ofu5AXhjUA6E8HnG++5HMw
tQEuYO3NJ+TkXzM4iPPfgu47SeJmzF9/UijRRnShwTG6U9hPB0EhBk2c6rryGwe1MzY3IvW4ukmF
ZNKi8xJWmdNRUR1eXWkW0fiBzFsAY5eq8qaDJD+go5EzgGSwxhqa7LznCylyItXADfZdVPLNnNmy
Mv3lWPYLJumTRW2z9XOi4oRTWiPSVVjPryJqaRICNsEEONoeB+X/zz6KuT5qFrNZPJPTm05rMP0X
m8ehKEInoYLfmGCb791ankIwju3YF9ReHagBP6i15DYgMTjg+5cuw+OujdOS4OA4m3uJv76NVNrh
tC2OAhYVe5sEQiGv30PXwHj1OWCBCA+o94Uw+BU890C4Y4dUkrIyGIm/uksVxyqOchFw2PxEpTku
EdHZZDQfR9sWrCssgH7t+3215plo3+Mxaih4zwdv6+RwpaoIINSp+T5a1OyH8Ok3pRIMIYdCl119
cSkgcp7pEsAoFHDVTZu6tdOXr6LQ+l1PxOPaBdozeb/2QmdAujcep16wLSqM86HpwAscxWYKKDTO
JAnkRHvXM63Vz+rdT3vvLyIxTT7VX0SoU3qsB9iTXJpxfiqf7OnVQ4q6/JRm6HLXadliniK0V/dv
A+TonW7cn9jEwwj8xtWvUI5HAZpcD2VPnN4Ew+9Usn75+JPlyjK/9r9f6CrJv18uCI5YXkYmnPeU
I45nZMJYkFxbN15fSc5aPXpo1NH88OjSfK65cQCjKXZBR4e7tOgFTMAPHbB5IBIgTTe8DiW2Mpct
dH1LQWmHZ1KpL1O/Z0buQGEJdykZpt6xTVYhD/INOISbM6nGSmXm2qelqBrUTI/WF11Ox3/8cD83
bA1uOhJAsimzGoPqt+woDAbMaPFFNMCLnULZNRTFg4V6Ii2tIoHN0Vzyh9jHaOkTJIAG1CaILyI+
F74U2c4qsyGjTKbwbu9LbbX9VWdcQFg490/wl9QLe3TQoKbKH5BcGf++hC12Nd5oOItsUBsqS4Ls
LMsGpJVkqlGhaCIYMl02mQSTmfuB4Kr2vVuz0z+ampB2uQyEU+ktouaYNI88COgx8C5af7c0H90p
HycUQwC3ZZQxolSYJZagI3bZStXO73RJKS/FfMBNQv5uqadQVDmjqTqcSiQOsm//NDL29dmnuue8
ReggIfrisRAo3xPQm/EgAadNZ3TbBWbvztKj/2bWr1QFylZw1RmKwiWVCzjmhjaLOfBmzYWrcxK7
K9fkESc+4mvmo5GicmdYpLS8AB64HRS2/hVKxVLSUSEvjUWTt77olMIQbNz75kr8cWqIi9lFfErD
OB7viRpCYXIonJ3gc4snSdnDKqoqjEcY9AsrN650+8RFuG9BcBuG+dRbbZGjHUPI3WOZsjsBi+mJ
O4I8ZmPud678v4URmaxWRNocJefZ6hvHa7/Vul0QsuzyxcEsQtD3aOwrZU8UyjIthreIg5mSg5N7
l5lMySzRBDWw0CCeenpYysys/sICpfgl5/5ZNaFH2bxvUQiKnzeg4mifba0KKBlnfTuQ8eJEDbdx
YrDN+YKNGRIihP3Q2EUHzrYKvk1dv/nKCj9xjLKl04PRY9HAxMu7i9/CUwwvubUhB86lDbW8j3aM
2XTFG4qhT0nQU+Q1Zr+60BEfKzQGSFIUCUaR3njb/M07dMpsWM18Z5fH/QN30XtRqnW5Uyp1IJvE
vOxEptI8RcmMbFfquk3vq+C8GhYVaVOKaFCnbTP97sRBYb30fZ8mtVHemMUVlXTh50nbX35jG25C
5rC0RWsTQGLqRyiXmjPXWh/7IC7R9j5+ZZEITTzMGnixEBE5C3clM9MMuHG/28GOD8gA2Nd8iv4G
WZPw5OR/hotzeEsNuNMzy+VuBI/a5Qko1n+rH/QXjuUOFin8IbSjXvwSuPbaX0G80SGduXdJVZ/0
cfRy+mqZDnRBWRixRjFk0+EnTY04P7HSvG/YdG6+x8URDMPH4HG5NFi7G68VIAkh+81TwaBb++l5
7uUDWcPJ8YluYtldM5w20MInsmAHOYzW91c0G5/v6pOI3wOylt9uNFzEL83whNmxKjp53H9QUgzf
LJWufkK9kDlvpeLadPuyGAW1qBmOn8+NaoEIViUFegSV9ymzBpnKAWcv84+ygcCFq8SsI85pYGrW
gsAGBjSXULdSCzEmPJpi6PMw7JYt3OdUX16msuRjjG+SwLzgdEleOlwRbjYahvUoxk9FQD27fHKH
1OY4TTsfebDI0Xme9syGM/B7zGONo+iC4OSm2hcBMVlDW7VrQX9B9SGDCac02sAs16bIDxIX0JCe
9MiYTU8HUBJkyYFw+gZUKb10MPi7gof/h5+8DBeosTPi5nu5qYLujIs29nUa8vxkmB2WHFmj68Eb
dEmm6A6SI4BiKOobqD7hj46rPdo2GhfY8O5EMUTtp0DAOoOPYORKaMKFETe4fzMrJiBaops+5x1c
oVdeO9q1Pdzt6d9HNTZgnKKuGAFY1Y7Dirvd2TN8GUTtTUmLPGUFelSify1+FO8LdHrqhkPePi17
swD2hWM/UAJcfSsq16H5SbRqDvLVTlfRIZ8umNXhdikoh4hwNUvCTU5V3eYjVfRzLp6Fq086ACwf
uQzAVMMstBFXNMXQHZvp5T/OD4f1JXbuFiKjB08mjbPtmiqiYZxK/vB+MLIm5J+MlMLEAQfpV50b
n2KlTMqmZlw3WaUQS9LwjcB/z8DUHNLWRpKM5rauqC4Ii8yLq+B0GiCETUaxCYtamYjvY51aWYRH
luDRGmhX3CrBbtpxQmxXpa7hm05Z3HQ8Td6906/obFNai38ifYN3bA0BjOzxIeMl66ZUv/OsS2N2
qfltNKfWE3CA3jhDCJ8clldZKqi8ur3VX6cYgWMRiCoSB42o5S0plyHQh0bFUH24lFSqaep0womA
HMgNAR7QwHwc6oNk13q1tpOmYgkGuJt03826rkLNZ/icH7+4y4g7Zo2Dq8P2TAKv2dYODAvR7+s6
7Y3QYHGoiVFVgOxC7KhUJhx2bN5XLrL/XhYNjO36rPYPA+5O+gdGc6ad3Vn2+n4b0b8x3GGLEBJn
VEW5BwaYxgNKSN6oBlN3ivrTltDHBq9adpsEBfh0Ghe0zjPceKc3ZcOxlQGxFEdI/egi5nRS+e+u
UlIScee3CyDraj8D3oLT71n3GuJ6dy1oA/hUBDU2j2knpEP3EtvQEx4bhzdE4Bd29m8egcP57Eka
3nRwbzM7v+s1EjoKO/JlCxzjAlDNkGkrfa4EBDP2IQuMwCv1k4ec8eHIGRTaGdZej/TH8FLFdk+8
NAQOSriTiuuG/AnNQXuROKpdwslEiTh2MZzO0fu/vVZnDeIg7xulPfizvVih+sSf7rbKlXNmpWad
IX6y7SJxqxKc7p6DUregHshAZ/Lu87o+3I2G/YJ64MdXrb3Kz5Q7ki50XI2lgX+s4Zhd8YrSiQZ1
LGD5ejyRiBP9LhGSAwbBwNcRT3kRO4V+I0u8RQsjEEbaozGxSTqSx2EWm5xB3hYMvYOb/2yRgOL0
jHMyLmu2/e5UpGatWHZdQ9MLBvKPxJ5OSxeVotpbdyrlReEy2Z4nxpXVwKkjntr7pFt0D+kI6eVh
on4hfmW45RMxukPZcDLzoQMBx7J2ROxKS4Sf7fEfel15GaxULpWWE8U6fk344cGnlip8c5WzgRFo
wMwi+NMI3SWsrzcDqTgmdkMMN7xhS/ynKHeVYMC+8YF/ClZ8HnDNgTqSncW0AAGeKIg+vYuykoOY
eNbpVExgSSSFzJXzGFHeDytVa/pvONtHB+y+gqb3Oyj3E3ST0owp6jTf37rrVxN+m1iMOnc7rxG6
dAQC5OI87/fvj1t4Q8PxxQimXHxeX3WPW5NdzjA0ZtOI1W4RkAOM7YFRISpuoF3gM5GTbLlINHlj
qSlQB4Euh5XJKcxw86Nh/Tm4Br3T/aTvIb5aVigOklpUfO/mkV3uOzV2eyKKVWll6C8ML3aDBb+Q
Xl5Xf4ar96emUVSkSYvzVG3CxIF0/ojL7B7Gih/BX5oVDRDweqjl2q7Ph2A++GIDTEh2rWTWkobi
5HiJGhRciEV8+fxqQ7B3OPD3zY3u+F8BDYj+HLfED2Q1kESIMPxJV1ez8il1LOtNvkdtP8F+foq7
+AqVMFLPs56KaKivQRXtM5DlH97/K+PhI3diFKyWuDJvWM9TsDeAAOMfTKmBo8Yfl+YkDUBih0sk
cKyntFrVxbHXc9hqGe/FbeyHWxUwiYduhs+JH+a7Iw0oWFr837OE4mOL/V2Z1B9hkyMJE+UZhg/h
2l0O/WxPVUQpGlpWwhf5eXbzheaoyAMGMMOazJy3lIEJZUncIHKk+EorPEHVk+5Wa3O8NRs9bdJJ
xjbctxn3k58hh8yAaKDcZncEnvYYOK7K/fL4+QyztqZd3wpaLiZHFVdrFLtWsKNABwGcscYfyu14
Uy+BUUp+HzTfg2lK7zbYlYsR8hViib0I1Qf+82k53v7YJp7mbsUG+YJbFaHDgjcOjQlE75cQj/aS
aRHEo9qCJ3S57+sMtFVb3dyRNOZMm3VxwhJbViBF//VQ6+H0F8LrJXlwEHF0BABAkahcm3d9l7Be
KUIqfX8sCDkcccSllosUgVlHb0nzQpCmNqy3hyayOHvnu+BxCwkhVTmiw9TCfQar6uXCxmWzpMEA
kw2mc+jq/4/JKoLOU7AeHTq1Vf4vtECNeht4oxmXzfR6797+XV++4mSl/LVTFTVoPyzTg9qLhYfg
hNtNuHAPCshNdsupxxGs3GO8PsKCXPMCvUk0pjnEmOAOHx7LW6ZQZSk2cB90sJ+76mg6r9hs90ns
5W2F+ZeRZerDk3us1egrxX+MmkQeoFzhxGxMURy/MHEEGNcPkO//xSjNKTJfSsfobWSjPWoOFVEK
CMT0lhzKFtokc5Gl+Pzzofnoj5tbYfoJne77i9Nem+SP+uwXqUXhWSnXlVq/pAWW4TuAu7yuAMyx
RvhVQGP1WzzDRJ2sJ0NZUrna8uKosZ/OvQ4OvhN5infP1kCXrYYYWwbqC8MMf5mEHlBp7/wlLvgS
5cYzhnTQ4FBoBkZn2Bjntkol+IGccuBrK3bnB42VE0Th/b5sr7ZyQo8b/B1jD6y1C6NYFzCrd1Vg
GVP40Pc8w+AFnv8CMp918EiOx6JsrjMRfd7tIXOW0Tk1MhI8RRRaMtClQwl7rY0CwfjMzLpDIpkA
CV15l5qMYbDqrqXvibF42vGSiXCmE+mtWLBSKJ+CJ0PtrGPK3DeU/EDJQwqQxCTvBx7vfCBZXgOE
I83vHuxQ0y4RCESMmA9SD3JCa5v/HTV/3eowppsQEifNpl6VE0ZIrr94XRpEYSxsxokiJ0SIvSBH
0zj3pVBT4Wgqy3NGiZcRTkF0hZhCR42AXYRuZMVjvMpbOR7ZNClIrqC7shdTJIPvAZtOM0+WndKR
Gj9+skoypJGQkV37PN/0MXq2EoOzQDzkCknEz22MgvdJwrWqWgnsNkHKE1JWDGmLvqYm8oV0mGZa
kuMVYwJVJkANG2ezlp2BLNJFLX7f7VJ5LhG3zkGZh/SiZIz4Xybt5q4KEiaVkgJaXKmAXpLC8fQd
3HJhRAaA8S2XbiGfRet91V/n9knDxIVseyhBhziUXxpeC0M6VKNr2zjekasip8VGISdjE/FwBlQk
VXEmD5SKlcHKA8Vt6eaxttThc4hlQtyOsKpgSDYPFKH4b3ZBtHg06+x5Jhp8ANduo7CtB+OgpNMm
3AD1aiFPfXkOIywltyj9YokLAboEtWpG8UhYGvhoivRzkxidN9JrmmnYPtZkR8JXeonPwijsLudt
cRp1L/sssBRmpz8JblhasOXQ81wf6x+8T7uXmINevJGakaVcRE6LxWd5GN3VFDtf/FKM/bCXMEIW
48QEDm6JRXldqgMBjNnauPypASqw3C/+I1wH+f9SaaZnDmpVKwly3q/rO5vxzDSvVvpcw1/jdaVD
xgvCLLmGjR6N94Ps7KLqUIwF/o0Yc5CEkxuxIf2jZYPgpfWnwoKDQVRIa3z/6dm7Qz+oUc0o8wS1
qG80PvFXY6ZVrnwcfO/52uDKEm4SY6kgfCMmDEGXIbej6kZ4N+R5Vzb+MZY4y+F+aBW4Sn1PyArC
VpTqTTkf13pW+T9X5laUHlGYprngz2EV1ZVMJOelRL5fwJaYDSHmUZRsLRVGuvi5cqrM0rfp4vEx
rT6hlrnCo/3Gw0L6J3Y+HlvqaexSNOA9Nye4H71qWIS0/W/dVkFqlMBNe+nrLxL1Q2pChBdemesa
/+azMf3O4WGbHReZjZRvolbnpUXE6RoLtiBluiYHrWSBbtUnZxEHvOrBn3rC6kA8I8SHCdQcU2f/
sfIqpMdVmciHx/bj6HbZJ7HrNkFrUldxPLwXfbmRsTaeKkKXpJnXG/YhNjPtEzDNRWqfPepGx49X
U8SoifZ01bcWkrr4Fn6nXJOYWqvJSPCg9CArYssTBbPjjICNzsLbS5V6DcYc39n8G4PB1M3Tgu6/
c+trSidDQVBaqRT338jTZhiOI6OquKrkozG1AyuzXZ841bJ36K/vJpRjhnDdwar7+YOnNRSGJGc+
UPicYPUO6NgVXFT60hB5dk/4w1oRahwfHAxdZ2BL03rdK2Zc9HQ47g8aO6kPdE6VYf2GZhqRzmdf
+vCBnGmsR1F6eAgVpP6ya5p03BPEOyC+32CQI/Fw32J7qH4Inl7IlPTc1R1PZZNp0XYy0ZDZvOIi
tj/pILLblEETWjyd3LqlUi/7eqb7aW6sHf52dLizOKsVAUBwvMzx0XgX0sziXpJZMSiVHl0VZ+s4
K8pYTICQCAQzA58pezGT6T1VwIeoNzJfyD7NdRkYjhYO+ERB6302Gdz2Z819PIfG+XJbcBIS/bVb
3UUuFVdL9GcUnE0Iq7kFpgGnkFWk3jiauSA4hbPkFHM8iI9L0kElk0VhpB1dlqU0MwmbCdr9ikCc
FjYGRvYsAhL1wWKUNR8cGlfq4qogVERbhN02A8OCV2RZ6SfuJutpBTo5+VjM/PmBwpkoCRxOI1VQ
oBaAbMnLmtR4GIUnCiTgAk316X6ZAOSn0FGnv+ZeZC3cm1q1TOdfXElc+undkoJSK6r/pQ0XVUw7
KBHhG3ta8DcD7PKUtQXj6g/PoLjJnFr974XDD6g7kA/ajUrEJlDGJebOZK+SIZRaNG8+6nNI1KnF
LnzafCunuQjOIE0pnbhkgYMzt4Eu5u6oWSn/B3eczTZalmNsJcbURhq6V+BkiClDspQOCkvoal0W
6GFcX6IgABu1qpavrsKzQde1CBRh3LviwhPYpbMPsWIuJRhH/g8SZ+YqftWwy/pqeoFzJG4J99ll
99hb+vqH1CI53JM4mzXqHlKJxsODs2mtBEq/F+fUA0yHtvLD7fPB8QPAGgdukoI8qnjw837jW3sQ
jegKY6tDZHqdH8wx5sZqFWLuulB0LT2AvaepybjXufPW5GZ8v4WanFSV827ZuZDAit6mcnX8yOtQ
JXqN6MFHPJF2ouleWvhD9LyEZiSQwNHRmc0Tn9/jvBhWyys+8pb6j9rgWjmcGny/3trDGl/+klxG
BvDquwz5DogJ7Exjnl7vj0Ofy/cV8TB2aZMUSZAMPChe9qSm4DknbJh0ND95IgsMsuJAEh6TpvP6
nwX6387rwb0Gwu/WYzGjVxcwhH73Ff4p0n6CCZnswGdxFrzjRPJ39FszJSsIRDf9woOowst/s0xd
3ZsYbsifCKNQ0uIAp0Frh8VsjfZn79ZJcAoPLIIls9aCv6E33NUxUEznI/6vV2ATSRP3rbxq3NHO
S8IW3mhByPE+B0mRO+ubYZRy1qop2U90WbF+MBHwT93M5iRdV3jlAUz4V/KNrsUDHv2i80iE1CUv
ddMPAQOGz04o1urtjYxH46VBBWcB24VyZLkA/Vf55yPqPxJURQ6cjkJ5SJ+syfzWsdtEeSa5ylYx
CHUZuYMueOvFldxbAKvO0PolRVdpqNbSc0elNjWSd2vuj+VvtCALtcov8FnHC4/ufPMR3mcbjhFS
I+w6qi6pU+FE1fjcaweq8AzHXpiDaOsfCaESegS/PvQ6AEYBs83SfJgscfFBHhvXzUSZnSocSJje
rA2zwT3Mwc/6tn/t/Oh5Bsg4JuHYX4q1n0M1K1h5hLvNO045rlEh0ojqiLR3GV2JSmM8VTrHt3/z
FZvqzZ1XaYEnL2OcuELzL0/xpu+84jBJCff+QFacBx+UeVhMmY37iWqhrBLQ7vfmDtoKI1bHui/n
uderuCgiBm1pqj3BfW59y9O/zzdFLJOg4538Cf7QNTL9Z6Yv0xXw74rMRkv0ug98EtqRzlaAbofa
JKh62mQx2nIYfhR3Iv6xHUUjQ6MlFhPuzUO1/l8ExR6morcJA+U6AgfkUUTA9z3/NnTRWqthnb92
bsDHVfjR8MYW7P2yCzdyWXhjQrm/04R5XML2baWz5txiegr1YKv4vVEJSJ0voy/UjWG2p7ZovgnL
ZrtTdaVFiI8rB0gKu1eaTh3TEY5E+kITrADxXIJ3K1bJIeXJc6MFoskoL8qMVS88/RG/zL+D4qcb
tmO1fQxAxtcZMwd0kI+Ev97H5vYldTISDSpfUjxBHXx1oX7Crv4XTkJOx/spiC0bSdO0xoDRidQl
6QRoQ8GY4Q/XtvkXmqyGAuXhDwD9oVedwFxRkIkZ5J6hv+ucKX7dE0x/DlB/mCDyt8aIKpQev+yf
DLV9jDhyh23vsAj8WMGxlcwuLoXlubNm7NZfWKMNDS4i3B+BUNHLoUPER9fifeAgV40Z3d0E6EiR
Mw9IgImQbtPLljI9+kbHMDqXSxGm0nn+vpvMu3Erd1A9JIPMiSQOYKjDdeN8Rmrhx/nX2uQAGeYN
Y5zLAi/4BVG5rqh8a4Icu3ttZVS4Oq0CI64fsSOaVQutV2GCqAxE4qhi0MLVYE8ELeaIbWSkved5
E+av+D3zeRyKWdLCvwXI+ko/nCigStD3GhPTR/7Ly77pj8Z2xWK1UvD3HItAfub/D0GjtpbizhmM
VJQBEOq10WOLwF4vK7yyIu+D/rn9s2oYufPINnNRxh+UzFPJrGBy8O41nAEmMFsSKVgEm624PGkf
0+HWDklsK6AD3VKOkAC4MulREbhwncB24X5KjLSbveCNmUv/ZTZ7P9HciORC376v4RdrvewrJS4h
+YrTVBYblfPRUGb19Z9z7TFB0k8B1TsnQvRk60nzIy2IuVoxIsqdxXcAvqLNpMOY+WxeQrHINc1K
YrR6ZuKK1cLWx6gVF9iVytn2gfMJxIB9m2/mQ7D/RURlfKYNUr6StD0nhOlVNolfkdSA2+F15l01
RySi61/MPghVbV473N0/pFRi+iV/e6KheLngZjM6QeBn+mWr7bpDWZ14V8sWNyayq0tA7QyEH/Li
MUqOxib7+6RJYHJ7HJoxfp6mwT9NPDS6FF8MmxEpIFoyEorFz9SeMAO4yMKwjlFTg2JPvjQN2OqV
zKcjVxDdxu2VpIhQr8goLO2JhNJeWNzaZHC9wOy3gdzJ5NQDbOE4EisBDYTVEUBte1p4GclZFkjS
PBeIzoZkTTYeNw2dFPhEJ3P85l6jDI8AFxtmYTuGXlr0AKCNOSkJnDP/WjakN6dv7cBZsvT9kHJI
xvTxI2KxgyHMVvdC79pL7Q9agZPUvDheR3CUiBu9AaQT4UXiKKyN3tu4SGp84zGh0NNBpi08NjVB
LER/b/cOuIHl5dK3MI09KRtUOddmWdAGYKKSGsN46C4VO1JabtY4VUSb7t26SMfB76wyNBW7RO8J
G77ABOh/l9csVZSQWVu3sRQB6/R/VqOpUpKOXxLhEkZW+RMBIQv5mc+k2fq9JjkVdwHg74GBesk4
YkPX5+9/mkKE62d5WfECPMxNbRLwzK84cPUhdHdfflJZ0HhiUyxCYjMI20ePrNFGxMx3z89K0pCS
pXQHYN65JAtrbnAv/3nLqSv3Q5ZThN3m68/NMRjrUAtf0NST/j0G04B2i97yGgxksRxQ1Pt4/O04
yE6JLx4DhDjyoH/eikqappoC2J6wUv/0+EuWqT1i9qj0EwNFfrcDB3HZARHAhgDrscd62181qojQ
xEfaq+yqKWSIw2zXHrFFfR07kXpj0AmFN009tiQkLiAXCPtU2eVKW4yzDp/zdUQTGP3r/JAcOI7A
+GKqJcV6UsLc67OiOhK1mKI5JA7V5dNmb5NP61pfbWf8qAyM6YUhQEJfJtxDpRX3xq/8R9vp/lq+
JlH/nXnzVMc7DqY6qPuxp6HqztsPAaihlSsi/ZBpV6ABLFZ4cT9WkJuLxKC9hdadTQ/eNR9KlYlO
sviQNdm0wPJT9/FNLlVfWIOjVZgAJ31Lccc2UFa25+pXDGG4AQnGpsB+HJ+MQqtP+1hky7ObqhwA
X/Qxq91oLMPtt8RtYqIQmZ6iQEApiSSfAD6YfTHxP0uIWeOdwOoNFN9PgCtwa4SYqHi18U5JD5Tv
0n++9h2zgMRaQXqtb+PnfNmApkKQb2xm8evMmgX43QqeWZQk3Y1cT4itHM+ytZCOB4TnE4aS8ea9
YW4LsunebFg4wK2Maq/KJNPKMwrLoFYeyZLWK37dyqFizWAp/mDd0nAF7YqGy8jN1Tm6bY+wZP+B
YZPk+GxYIGQXBSTQFcwImb7piVXCNwM3Jg+PfyDAxbzBXBJ/nh93xp4jbhLeGNPX/Zo0cVIrRWCL
nqXU3NuCj2P4P1WQglrZvtOttNJulVQ3I2jF/t79IgmLB8NNlqUCMxvgktzoYdlwkywPuuHsNzZA
dQq1t1DRwmzp/V9EUTQvC9t0EtpcPG/vqkmL5y9g3JCcVToCubiUQ1o2cv5qmUEKyph6uDU9Kx+A
8F6K6vegQbhFv9laylMwCjzfqZ56yBkRVQ8ERO9/9wJ/SfWcib7mfmnR/sqsT3yZ0Eg6awoLJDDo
rIxPnGLdCKwHuXIvhvDR0+QVZuwYBZKXBOsQ+8qR55i7e2OBXGFxb4Yu+UVMVZ+KyBT+5FJkPwYF
bC0+fjuOuQunCrzemlxxJ49ubj9Eysp3myopJn1dxG1SHuLpFbLc6gdMUiMiHd7+1pcU0bMPngEk
qZZd9RpHPhLNVPBLIHNk6CcuAIG0qtRJp06hoQkRDcfbZDNXcua+J8h5agtzfnu6fA55IbCIKVSv
8a8yylYNnMLtF7NXzuz7P+87eHZ1mD/o8+ZNUdfKYA0nV4h3Qgp22hX5nBl5jXlZAc0YNJ/iFTJy
YCkNf8C/VwnWaVOVSJuMZyTh0gtoXWeh52FNEgoL/1l/r1wpv6aUbATxlPOnK4oyVdsKFFDEt6/A
cyQ7Fg4rjhy9PY1f6Pik/HiAIDcWsr8o+tDoZ3l18iWRXrBKoTksyn6k4tCbf+Zr+Fh59ajv4j2V
6MB86wz2nb/9hi2btsNow0QtGfwEoKlOSCrbeGuSffLNuwqXzC9vexTlzAeptOqGpKd8J4Tvu7xl
gXDx5GqUeK9N134lsaCcd69043Pwec7Q0jZwTUhHzf722wKuBPcE/nFXizlh8shRgRAK2xkHRKRn
RHtXqowN5PiH/iY+ngfjjZbc7OLW5AItm5zNxCKmDOnS6QlF+swFYrmutohrdnezAFTUvEYYFt3t
Hn1qpCjCeHSzv9JXQ2vRUagOH2ChwjHyLNnOFipoCYSuWG+Rn0RIdXp2l77iaC4FlaBBZpCo6maK
NkTpyVDzoj8QslQVlOM4uleqGG/mkNcbxVHy2bReYxYpCGEwUmzOA45iilF3Gr9Q9zm43ZwuS4+7
J2x/NdwAyFE7DDYfX48IFyuMGJ9nzy3hzfMN0ZA3nd92aLOfsvxCaoEor+2FUuYlza0gf7yFurWt
rLtPQZ3Uf5o6u4QRZQwd5uB6Ee58mRTp0Fo/MwFt08Vqw9+mrSyKXlNmTJ9re9ovcyptm3eY0BB3
m1IhCzWc1FwN8TZlHFvZYIvpaxiqOE11PgeqZkcrKsjM11xLU3x4n+VP5N+VEJOeRaWjPCUBIJLk
tgBOtQvjJQ4A02k2Xd/8XKxuz1Zm2UPvzNV6F+SoMVeVa3EsbOQpbEU6UK5NmKwtcCyRTUZACPxM
EoR3BtWkgNhr99BxTZkKTLlKdg6kSKFH7PTBbYBAK76UAz+aznntBEVzbP/lw6PlRKyzIIrewbhb
yLQvv+CLV3K6KJw8ZyZQRlEYS9uPyPDkkS1/Wut9F5TtA7NGmxjiWMYC1/deg4oKmnxrCAnA/OhE
35ClbqrH1Vs9RJNGgqsQn+yAcjcNmzLPjl98EmcGIFlfZFxKYfsd7O7tlS9Xb9qS+eXhG0RRhUyk
xMHZQ7NiGPJpJZlm3QQ9T/I0buOkcWpN3ZM/lZ3icznOfloxLwtC3608DR8/djYCfmVjgae6Ho5e
YVu90F/CrLtknQWOv4kFiNjvppXT+u3HBEvO5VCOiE/Ylm/C3RCpBgICQmzMS/iXU28idbeigP9q
cwshJnshvFkBp4QbMpQtTf+Rxq7ZlkBI8dDzwE1x2QK8OfN19aXaW1wyR94RWfKMtVULhUV0SQHB
LuUm2hyp2V2/9HmyjcSI/pV14QEQC821Jr/bEmdISLhUzHKBvOWBqGL6z3v7FOcoAwAAdbiN/7wq
S3SfQ+773N/Y10eGqabx08KxYotj6M9f1pL9eg6shM0mma633ceQvkwIvsHnVSDTkM4BNH9I35/d
PJvRQdyFk2GwK3NSzs0bFB9bIf3WF+3RHcnD06xZPalngKVok+KNHZ8lkzswaHpgB2rJdYhwt2AU
z6NVTWmjumAfR4PpkAPthl1PZka8X8jKjROF/UkB5P3sqrsC6FfTXZomcKlSYDXdb9GOSrUFPwkA
BVQb8OPta7PklAiN6K+XIQWa9WXlIEnjugYWVzDxS5oIiI4pKqA1AEKHUzRmDt+WmQgUBBIjXPs9
sMlS/XU78wHt7bJoYN3DgfUEd1/7Ycaj2qQfyUQlLr5xyxij6JsHnOtUmPwJvffZLkv/q1Fsx/IL
BANDeM9fL0uP/GOZGMquH2L6PKItFfC9iiEnj9HFPmA5aYfvUOmUvLOmlJvE94p2ptB/aJAhEHY5
tfEN+ViYzP6FtzKYvZiPdZ8JIGdNxZOhTFwy3FoWGaLobV7TkH3B4ron3pj+66+s39eL8+Adl6t3
6M3kzh+xjtPUFzIEO4naQl/BPPK91bMljYdzLkS5KMBnS4eZkFJK08XV7d7Q2R0WQ3Cbb2b+RS1e
McrKxK7VyMmOtRhMAPEEtIHUUO1xiWaQa/xLf8HNUUwA1SOdjDcJ2o18KrO6dO8Pqtqqogyo05bd
uKaL8KQWuCnqVid58u/0dnUrsqADwoo5Y9SzYDceDB+NQuQqG/UfFvPqMqG3VQcbBiC7D0Dc8YnV
CFVkf2kDvxcPelf7dF+4uXWXlLTudk5Tb3YmHzJ/84mJfUVK4fqj/dGZnyjFQCHkY1IYFLD3QWQj
WruEXTaFRSzi3ePOKLMqlvFC5sD5hgv0zknR0Mn9AQmNn+Md6UF+WrQBm8WX4jr59mcBbZjJ/S15
ZkJhDr2YBkDeawo58RMfYiwcUwgGtRAiUHvNN2Nz+lPxwdNzU1lrMLqw/paH8WL+/KRHKBg+Dkaq
BCOOcMESu4JfV5FLK62bnRo3trI2Ird7T155zPGgFlaWR6dNjevxTUVN8VDPI8NUxgV9Nna7So5Q
lVD1YPyqtJ/Fkl7MF2lk0kStuSiZgCRZzOVASM2s86HtOLBpXA/NvDx4YPAkyXLt64kO9OPlyOSO
mzNVO/C57T1OEXeQliTI/IK5n4Sf3jw30FVM9KHqWlsFxHIeLcqYsX39wUBWC1HCjIvy3roJeS9M
NZBHdHh09LR1E6rnc/caPScrT8ev4d7qGNv9pw6LuVTKA6igxXf/DMv1PNOLSz2Rzk4dhlYEd8wi
0Tun/32yZeZYGdcws/UPMRR/fK6koSjesPreLuqM6/HNFPzxjQBrup/9WyGMeowc1wtZjEPxC35S
HZ2MLBYD2hV1oYL63Xc7tQJje/h3FY0xWhLxTKIqe3tvb1BsCllBIPIpayJ5q5jR0+41VSbmtz2/
Huy+VNzllW8kulkTOhy5G8A7xpfvALKQFoRtGEARxJbrKf7GAZzoBX51Lu0OhWJHIQ30SSMo7GMV
i0KDacN2cQ/GcUA3hfMPjVzt9NMVVi005MxI1WvGsLH9I8wrDOPXPALcE3toxDyHMT2pmZYEgvaf
S81mF98kyI9xWYe/4F12pAOAzSaA/y+GpT6eFecc+Qsn/Kprq6MX7NlOER6tDMxXhQoyvRvTbei8
hPxWmqBvV51LSgwqUTsoZhfVfY004vQG1C8I4gXNO4MpAaD5c4G/bbhANhN+Pv4pZW1bXbvvIjks
SooeV2a1/WuuD30eHWAA756oJKagSmviOz6bq+PCnyzz25BnUyFmh0pxeFbk1KMYlUvvnHHJZJ5O
l2ur8lSR4UfvXs4QZ0KM+h6O8KelCBxokrz+dbrDUXAP6GX8xyqmZWnljr1H5+3inApP0slBrpzo
MNqHGPr26NauoSh5kdpy4sf6hIvmyIRPr3aKraCMS56eKex/OKclkJtNKxik/rW4iQpmdOrWPA7r
Ns0ihwVa23eM0IehhFi8CnGU3AM9IBZmv5T/slY65i5ROC0X5lQ7sDX1EPWq/ZElFHoKyNcymhKF
gtRvaZ14qaaUjAhmsVE73IORCElNEvi/Hj8gESxdL2En5NtgN/Py/4LP8nPrvub2w+9cSwS0tKge
YbJlLTawJBIIqtS2bCh70xLSWLQv4Cw1KKlmpjY32r+2QeQS8CtKE8Hvh1VJ0lulfvs046rNej4d
67orwSk6MrkaNa1V8mAx9worhT+Xyo4brJv0HZgjn9iizSaRq+CqCKy1bwcMEvERwQjpgxh6a38j
8hLHUwZDnNKaAvH4LEuDYRFr9E1gTW0M/+ef2E6eJiW4/edsdnNVb6uzPKZUYxyPNUF6bwuGEa8i
ubdxsEpFwJKag7wVMFActIT0nVPxqpR5AAay8rrsVErQ/rEHh0Kdkk2gI4VkKam4S8q5KqdmKHwh
swzEDVI23zXEPXuyymix+9hYjIWa41OlYFfglZwa4lhW17osHAs4+VULkSNGRQ0+bTuDch15nA+8
YsAxsc5gRnFSsnDm+nd5J546bA6XcVkT5hXAEiX1HpRzrjfUcRYNr+sQ8D++W4tvsnFNmcbChWhb
9IT38HGpCF74XNNc8dfgAy2oaIf0U+XlihKYSRPbUetNgaNeIjJJMkQMVkh4qrZif/GqTchjIRGt
ti6chWh8vuVcHcL2kI9yATw1J9beTF1VuJ9h+ASFBmjqdC/1PhRxyEiITz1HgizYx38AJPUiu1wv
UR6eM1+9TlYA8A/4ZVzAkaLy251uqpOuDpSSBxhbQvCFjOJ1I82y1tMNL2X89Lhf9N/tzoMjb3rZ
hyFNQihHfEaYpCFt+wuTisr+mw8fdqHcNtqm9YHVKtGrjRUtrJU+uvHnVPr8sEofncoGE76DOqwZ
HMZYcgNZLrfpFie4NtWTA3JCRjd4jbd0Tjq/ANUQ/t+QJbr6JRGpG4EBcYr8E4zXYl473UAQWW3b
D34KEnckaV5ejceFhgzm6hIIQ0z926GptQh1NLpUE1TuBkwXJ7d/G4YkkPSZmnhANLaScKqFGAeM
q/jvJd1efYJ/4vg1aSJ7dVDTp4EntLX6O/vB8SvWTaPwTsxqcd7nJU74UfnqGUsN+ffPWa31yTjR
zSf8x3XU/ttSs5qzOzjJ0I5RBPcZdSu8tZZcgpJOLtKOWUY9EqoNipNiKXwt6K44YTDfdJ8zUXu7
XRayVng/t0bbHEeUlcapr45lYOb3+1WWpKa8iejr9wqXGPHFJNqoDSl0IzpsxpDPqY5SO+og7CUF
jKslyrl2drg904ouphhsr2jpo+BzAgCBL/uf5M2UUvsbSNJ4mDdjZHAc5THkuvGnTsTArC5RCxjq
hdO3qbkFcyrn3JL37fj9wsUB+lgZH7VcqGc8xtDRGd3qspKrj3PJ47x0RIHh9Hvw+1ie9RIXTSJ6
l4bdMLleRr4zicoflqYoLi/8PwdhEZ6eG5b5s8Op3H7nLpAxs3HxQQ0lpyfe0d6MfaLGd3mUag8l
vi0ZCF6p8Rek6gX0WaH09g7AW7UO59NErWxEy4ZwrDWGiWyoKEFnPAB27//NL+8wCdZeDe3oHe6B
sCLyXz5XVHSypGlg2qCGYy/jgQ8v2Q73rJMIyp9GOieTLQGn5CtWJG5rNbdzb0x6NSueMQmYMkDb
IGX99h9Mt+SPH+Q29EspbBRU0BYCpKxEymkHbLg+ZsqoN5MF9pU/itf/IyFQTyE41JibIG61KthH
YKq//QL5+8hq1Ai/ZbgjdrWhNg++usdW7rce5Z9Urx1epZ1SZvbQ26VQZDt5wzn1FqxUttUWXomk
YZ4ANMqWtBmwaESBbGPVeDcTxFlWUX/VMvCgTMXEcwXgHUp1utnpI1mQZciMTDmBnoatThoOysgw
0J9yd8apv2LLt+uuyy26GjJMvZm6yfmBF5OyISkQVvHkkPBT+1ryqiJ/j8KpTZ1H5MB8A8evS0Rb
SR6K0O5dzf5xsarTDxsAgFxd0bP+/r8+RLCnA2zpQHR7nNUI830J+GLHKCuZJG+MsndJ6w/kxoEU
Zexi2KggQEkb8e1JFLyysWmgMWk1F6we+uUmgGClw2aamEmyVKzqlEjWoZVpxC2Z8XvYwaNUpSDY
Gm8r8TYgkU/Ijp1w4sOo+NQhNUrPI2sBM5h9QBBhDnkgvOq7prZc1BgC3SAfsc+KrZYMwE/B+X1G
a9zkvczUFqumwVtrUPP948qz9D2yj2w+HeML0/PYqlX46qUlV24KEVm1aeHCl2gY9Dl9g8A2S9RM
0b9rsDE9MBqRmbkaAmWqOlhq7/rupzRoT4ppMXec+ArJf1q7jSCmAJWo9vsipJAeUbXzytuAUu2J
HOM+wGH9ShgGyTfHtH0yrQg+qullayOB/6VaHRL4bPIXOtBCGl1eq9fwCuhKdoqVBI+0Kl8S53cG
S/qd21PFHllRW/GEDrRwbee93YJX1FkWJrZC9fUh5jhGQHYJ1DIcD9J1aOPH06feJm9NYLQEBqVY
Pyol4C8eGMQ/viitZj3lITdj03aVrYh5qgW5ZYzJo2+cIcZj+82MVVV+hwuaRlzoY6aY9f1kB18N
4wVN6mxvxIGHGczhP3j58Pvl9oMGwiAQeUL4dYFiIVNAKtEVAUBRpxg0LNO/p6l0wcxqAggTq9AD
sRf3xxDS8IHVtY1PU2whrUJaS/t0zbR8GhX42Ol5hgnbevNg0zvVb79efBjlVmMS59CfmOkD3M7Q
EW2Yz+VZQQ45FmQOwtCdY7/pAvkaAE1eyfirxB1QBQB22BDni+/CAin1MlaXWzdMQCzwOqn8c8X5
GLaDcxQpWd5W+qtr8a5FxMnbH5fb+6Kju6tY0WnOqH7pKo3nvEkCn1l2KVB3D3VVBm4aS4etMIDj
Lv+MXLqcmDWiji+djM3qbN81bP86p0h9JnaSBI2NLpvhkbbvIcsa93bVs1nzsT/z/5A4DtEPJ/ew
jJxLZXbEhKqNTisJnMFtiY6sDU7Ovub1YwwR+99dYOhpjEGfCKRJc8Z0sIGJhl4EwWfaO11Vvbjs
KHlTZdZ2pK2I5XXqw6dBjb8dQ/+IZMiwgiyVWBfc0z8YKVGV2YRJ5f/pGa5sahzUnxMS3hxjEcSn
V2uFejMWzXwMd7r4zDOVe93FKB+BX0z+y2l1ks0e1oIviVq27sdsJiCwGCPZWJQRDVdeos+NdAaX
RX9gAATPCv5c4KwID0oDn5aB5qxempbDGSNYw0xXWN2IYSrYYjm10D9NvWBbuscJ3p6KomNAjNVS
HyWOLYbQq261wXMHUCa1IthljMcIturokqAnmGeRqCd7i74Gb/lPIK5Mqjqtc2YMKA0fpH2s429n
OehqG+JPXyTlo69Vp45gJZZDWh4ehWBQp9Q5u8rc3FaGl1AOOgQrHS3GdSKo4aW06nr020FmLAtZ
JtVtah8aGEcVmYTnTljtOgxHFvQbZ6n/tkLYha4GCWdOQCA7cpU+OsHbNEM+L5PLdotr57ZzKQoD
hcK25J38705n8KjO7iQV5h12yR4MtjFBsy0DRtWltyrA0V1k1wX/NLm5ikbzdI6bTJ+xY/Y6cDRM
oEQGFS6NUtFrpSO0/tQ6kHHKDWAAQo2Spy16gAkBI8akCsKF9+O1tG2Cwgvf9mtXwhJrf5wRSfj0
46SSdm330MyxPmyNR8YM1w4HBCzNZVePv5qTK3NDki5d+Gc1914QfDauGJrN48nE2+gq8jlx4jce
1N6mVkR83gpsPT0h+GkvwNrIcENAzmq1vR84kt5BUx4Bfll/y5ms8CIPQvQgKqiwSFG7vpuE4BEr
fJ3E0RbLS6uOtewc/+lre64eRyIfhOOFIeQERoX5xDyAt0/Ot95RZCMyPmBnXEIlSSek2B70sqGz
ifs2FBcHZ8IUhmkPOYZV0mPumNJ9CQLOoSmGUElHDCpLpI/AsLt4IT8bPAWDMOubjohS+N+kXnFt
jDsBvoTcYCHXjYnzDlgsvQYvkxfObKuCCx92b10BeqtuNvqG2rGcgDk4oFSdGjiCJ1sJUpBCYism
++j1QQ8oS7qBplR73in/zda0izJF6jS8QAbug5HUHFpKb2E9+THjqOQ2WEZKQYw7pk7d+xzJQru/
aaaAxPhz4eAwzY0CKY6fuxdk4/Ac1+U+VbZgRIcJYHpTigwTmyvaprxBxo9zhCqocEMTFLWvziV/
6+vJcEGoFYw+KJQiHDpEp0cpwIa/j2gF9OAfYXTyB3sEHhjJg781Yfy+M+Fi/sQgWqjq9u9dsIOn
sESr22RiceWZL7Vy3GXQ+gADPKKqdEhpkHrOb4QjXKzFJV2hELuWvJdZRdqpatv+xz7Tnl/GaZ/I
QsT4r+6k0OG7j5JqZa4KK5uE5aNaFMSe+UI/p7Kqt1zw/1UB1zamzbepwbrAvnl7OURu2o4jfS4+
DUU1AwpsJ9VgJokWzKgKSAnIISk6XH9pkNUH1oSYkP2aUjNwC444Rsrr7y05VKlDfrRPAAjXJwBf
ygZc4eHIUgq36YYSx1ruuiG4P7o7RPz/y6Qxs1mSCN6EFM5FwBQoyim/tu/H/HQalJXB2Qj5jAZ1
BTMryZOHsBy0M/K5Kt3YryWYaRLw4zeb1a83NI8qO833Uw/UlUeLee9R83n9ImtZeZIghAhIaNI5
czP0X98KDDv79feaWu77LS8T5ujIU5dbhQ0b1+No6yCVvaJwvNf5F2UdHywoVyAMkawMqkr41zaV
UO9E+KF5PypgK3mD6Wcnszo7dw8uG2oy1kxSbyvxv1IDz3j3K33sf69Mfm8UA6e9O4RZg5EAX5Yc
Q318fOs0YcHUl9y83u91kk04kqDdINSS7/op7TMZXbH7xeHTDVww5ZQWhKjfX8SwjILYEBBJrR7z
WfT2c4iVLRvZfs61BlEVNy/xjqn9UgeiB2qvnVwmtjUZHzNWxp55x0IKG10cm/4IwidKVRVlXSIV
YrcII8ENFnpAmGQNribwZ0q0dpcLHRu02Xev7+Q1Ec178mgauQNnq0Xfjil4mU/5i9ibUI1iBKme
3lTX8H4M8sEP0ny28nfg/gC9Fel4QeV0tEWIBTIaV8b6SSHpJpyuvMTAZDDnRo7FICBhzbTS9J4W
/OPEgKIbZiqGpIvGdlaSczATmG5EedUqIE9GBdT0kH3rOEh1NmL/642YyBPfzkDghcIf7q/UWds3
GWDN1m/uqH3E7IYmlI6D+de73xn2y7SHGjNTIA+BwK+xPeqRc3sp5umBAHrYCLff9WNOMDw+qXH4
mQRlI87GWg+QC9ZjL8mjhxUoV3R9yshqx5U4TCKTrCaHziOeHQ+NFi9Zi2XyO70SMKrlgoSaYxC2
Amv5ZQ9AtZ8OSovR5DlMPKX7v+ll9y81GeF8w8jep5438udmMpdCWBlvV3lEj2eBtyuQlf99US6u
rdy0QWdHnBQMN4qF4AwG/rxizzicCR47IMPun/an7msBw0QlOycAdnkD+1SlhcdxyjvYFVCFJ7m5
k06f7ro/4uw6iAesqc3rYzZlvP3MJzu5d8pflE4L7+cmtLK3mZsGX5a0Ch0zXD8+GtsqtbLxkX6H
+z86eWnIO1rBOnhshzoZ5iXkoTwyxsUi3ICuG+bG31lnS5/UH5R/uA6icy1VIuFf52NSxVXc44Rq
KxI/Bb9ZOBxRBZpiQ1VhjlRt8wYgIjpUN4HDcdTfucXnx4zM8XBxvqwbIGpwtZ0fRj0nlyPi0u7i
3smKsDKaMiFP2zrfJu0eoB5SzVIDItLM70fSWUWXnnWfBQkdk+7WrqJAnNGDzUUfJUC4FIyRcrYM
fvFTYiOECdbq3OXzaMlPL1nsJijrgwAJaJ0QdB0lOhBn5OT0fbV8Zb2Bf2S6gzhfSvMeLZff1t/T
lED1W/iv3sDFY2h0zHooY8ZBH1EvvSgx+8FVDDPb/dZH1ayPUdInDo2vfsH5joIVGmkZQuZiWDpz
uET6Wwcdqbe3/H2iGh3ainFLBrrG8JvItAp8XMtoAL3aVOgEKZLYHuVdk5dH1cdBEk+c/ncwhHDs
G13rZgkvhM+psxqcLSYq8J2Wb99vk/hR/LUtVUhy6+G2DioBoaAxDhdMh1EDdmxCAn3NyTjkdVFC
1aQ9DLz//07wlhXAb1LfhKyGET4LIuI2xJPJlM8qNR9j+2/zpPIazrWuXDGku9tiZxvXLc5o2G6N
Gs7CcN2/iPZehWUKIrmztR6Lg/38VQmkl304MHYzfoznzxOjtOuXfKa3hU6ECaRvFsCnCiLhKh//
ZFKnVNcQsMZZtqUqlEpcuH+iUBywj3g4GIWeUe2W68/Bjn08Z+lvFrDsxOdkAZM6AAZs+qbQWcQ+
qFGmDPk0v9F5IljVR+79LZQJVD+FOaeVaAXLB8IIZq/X3Ls76pHsncf1FQcv9Wtah5LKmnZ/5RGZ
rjvWvsEdIeLeGKRecd5SuoFMarZsKOUNkQERE/WuY4QoTKtV4DfXz076C2xEgcxpaHxf6Nwa92kW
EWoYR27d4UTDDW0cM3GVbVhCldvL2hG+ikeFF8lFReiXOXRaC1lM2PlfPRUtvSK6Y52CUx8L3vHX
4LHwgyJrtFpJquaBUA0OvM9XPOdzey7JuGGQyzR55reL59H9Lkic+yr7pZ8Ts5+leoK56wohjKm0
G29aXn7x7cpqhwjocri9R/yi4U2Z5Uh8JDI+6AIFyk9sfandVsZ2ucASJmfcghAQKZwHPYdWH2Ex
aBOrcv64OE/u19wP0MFBYp7MjdktRZJojqodeCazu4XPUjulYVrxcWn+cA0fjkePgz6I1JZ/OLUr
1K355P3OdNZ2IA+3UV17b6gLfid7IlCD85hDHbtBb9m6YdG6+kZbWPg9TK6tE6ScirhkffMWqQUs
erhM8hooy2HBEMm7W5Z3tgaCEZR3yZYIUgwlIUWJQDx7CkiGetfXVvUwBj8p4BJBTo2Z1Xa9Um8X
S77uKr8RgQWiJWbPQ9QbNLU+QzgEQL4COOKuXMM8mn2CtzglMKuSyXUBPLLfifDyGf+JGXJAaJhU
FOY969UqNi+ZGXQ17yG/3JaHFq+BIChz3jE94z6Kvv+0quymCHc4U+EO/JGBjLznzucxhw3L/jgq
ud3UYkeb1mBgQ0qatLDTqp/GjudJ6788Lr74dJXOHF8uDrwEdjSE9Uo1gAJRuZ3aVuE9c/Dt8Tc8
6nfJLvkkd0xVz4cs2K9p9Q1zV7ay3jBdSGgmSL3P2z891cje+mwSEPIl2jgp6hjDI4shj8GkLxRO
psfwE9YHj9Mjdm2SrRze3NPwRepv+rpE/mpNrkm6Vr/2VZ9AuMAYbxa1jx66uLrQqP1ExOwq4Xvt
FwPgUMXCdKVgouvzqYOC6bX/rO8H+F7f2oPGlxb4XPPh+OnwMU1AaV4sbRrdTX2359B9JU+tNgQt
H5l3WtniYHSqrEnBNfU/OXbd8BnK/dOcSiehwHAF+jZ73ekJfUiPolsag6bLc4vL9AAoOV/N29Yg
aOIASwE3pC9gnAhg3wGzxlC7yyfbnzJmURyQdEok8JBxDhEHxw7CSyGfuXZqhkNfDmGDPTFYEH6T
IN2d9ZmB1pfwAT124I8a9H+iWZmdBVnJg80S0jZBbmFHIYNSqBQvOLRQVP83pvk2dCwI5FjQG4Ov
Iaod0uwQ4+4aRpOM706q6+hdV0cdNtBm9qnaty1weilsrgsoIu8VRoR2UH5oDkv1jXZUUkYe5wtx
Mds1ofxNO8DmdXXKa1w4T3qinGmcpcj3Puo/PP14gFsRqcGUidgMsjUxkiBghhTygUZVjNn5HQP+
vvYkVcOFjr7ShYURTI08bI4iKN/d5FwnrePieVJDBRUHWfoq0t3u7SpQhtPNcVhc8PAZTjM5b80O
ZCphwmOnahEVBKm3834K+rHxGDRQwHxIK/DGT94EdhoIvKhNeDXDD/o8G5LwJk0miPs7rD1W9hTm
mdZhXPjpccCF7j8vxjs1VCzGza8bN89S1drgLDIXSST+ngCfqvXdWLywlwlZVSaOKnqfNiDESePO
wmLnOaRgZ/GJoxOZJlT1uinCTBuQ/bH8riAoaIzXawd7BXaxuFbaqrhEMvi60EPidfDmWt6DFzKX
hGi0CUxXw0AjKMLBt1rK0Agu5ZXUzKEpwEQSCFCG62j/bqMZUffSi90ROiVfeJ3GKQkYjYkesypQ
cxcEvBhsBQiJc6BIMWTl+UNVrNLrG9hvt8Qv72Annhb7itwHnEHvSZ24gmO5cYxkPLWN6u18pGsm
Q+obtZ1TKJzMad+iJOhWl5keeIxSZxyD9CPkXAEN0BBQMizsGmecFiNnpaa7bf7yrOsuxV+hdokq
U4L6gJ3Fy8TAl7ZXMDLbHKEZ82/QXGd0ngO9Sbyq9OYV4vybI8c8NA9RYJF1kE1qMqOjujVs/zhC
XkhqPauHs368L0NJO02TmdkrjVxSljXb7yJ/bvDj7nk+EeDOl1I13GkSg22qNOPoeRgNJdgIZ4gw
1rIjp7pbVUG8b3vGevesUu/P/u39NIoSrYpWwe0us6ClcsTx3/7InQydtI6LSqi/7CP8FsQcKbZn
IbTjoujcWdlQy7kDZbdMClYU9ZYB6NLn1d1EHBEyQjiiZZzPNrQaja9vBjYgD9T89eyOci1X8tfZ
uP4jSPtoMLIASyxWx4P6cxwEXljtCoAxjOeEXjDqCRagm62Y0JUvacHIEDoTtNKtSx7uiO9aq3ha
FlK/ffmR5ih9jSCfwiaOZB8U+0vezIsZCcroAhP68SFk/zMJHim0loIdX8bviFfWBDfsRQMguq19
VDqKncClg1/DoEssFVsqFn2ybtHxkdChW8JdGZFBgn4wt83BnVOjkfzV/GpvLMf1g8b8nB9FW7PM
/cFD9rU61MTThE4P8baokCsiTlkqlUeuawt8bLx1Af/3IMomUQPw7Yu7BQj8Gv5rR9zT2w8lJ2wP
HA19S/X4OQK2akzcwTsfEXcwymLXCaI8lzUbhhk18V4i6q+MQIvHqarWI+bUvUSbY0/3dTP2BpDc
AZ8cepqCf4PfxIUuK3xYG5OwHUZOoVirZJiG97A6qAr5kZLzfDXEQcXSRPmXYl7rb6V/urmAYbHS
PlDOI8zaMA+wotR18o5tBTN0VpvgAAB6H+NF85TdxbVQGJeg/L6ix0C37ZHP9liTvWH4KAWNz90P
11DSMOS0CK6LRLFAOf66a6QOv2W606aPulQaEpEbo7IopICseI8wbs3+/imRM6/fT1bs43uumbGP
kr4wsILGQzLrFENIoFPRXfpuSyH+xv2GTqaytPfkvpi+7dWv2yVjnmhKykUws3TrvfrPF5Fijkwt
G1druM8XOZjf+oCTj4aue9bFSDhnQUXSBZ90kU9OMirQg/qwFh/mQA8wCmUEShyoQT5Epp2ok6/s
YGpVJ+Fq2SbH0/6a5oRYwvEU5NlHckHpM65FwhbpKRkqy2j4fhORgtsip1M+muMxT5s5O02cXpqH
c2D7lswDPhTJ/7k313XhLXdnDO4NhhVnl5j5iTrGL4dR3Wc9KIL9ePuWcon5BFkBXtVzhhLRXo4m
FcErDVzzgj9xamnEIuYfd1TUmvJpfIIbloU0q2pj0nMHEk0pB32GEpTufhBtOBs/wCNVFh4momDv
BKMdTptgyjFI33bL92iLxno3RG7pCOfTL591f51YwydUvIP4+pImMqXboK7viyU5SeSGqb70KEt1
wd0FXg22f2bkw96uiVsIrauFBUiYb0e0Z+fAKDYZDJLOvWYJWCY2apeq9awUQXUVqNNjTTY4mkfD
TS4v4mgZvKzd6Uw+XNOTG8NVtsexV9rJBtdvyMjmGBt6Jhmk2XqAXhqaV4XNSWtyPFZ9lnWvoaUR
P1J0gw2c+8PqH5iHkEd0bZEk2AEeXveb9hN7dCRC1g477CRcPGlMVXxwnNXJ13NW9+/LAQ+QYh9E
oyKlUiuHlCkL0Pr0uf5Gcg+NQMvJSdY8sHQs5x6dDBVS+dYXwISU4yZi1+iU8xF7q09q/MJpmxU1
Iz7o4hgpjGLw8IY2TSVslEvhWPECTC8R3uk6gf28aOEG1YsTWOv334H1sMS8DGj1oMPaEgmTogp4
3iKNnTy+VnXxMdmIJDAk84JBDUxoBz2xBB7WSzns1AtVKVYCQteuPWn1c7FuJ+mUJ0fBjqazDSrQ
m1FJbkNB5nwmP694T/nzxgg91Ll7F+QoW+iOUVEWYpqUIml2Nswn1i7penFvx9WjNZK6tnR7MvGk
UtlfvJ0pNSndWkuKVz2Sm3u/czGuok9ldj0ERJKCtnjuKxbyGjINEHByEtU7C0uRbULwHCw1kbmk
0gsQr+EE21IDSyeVAeT2/7m4JzZQepXu7chB+KywwKiG6j6hCWMH3r8simA/gEom3YwXnHQ1ujT9
G3dwi2jjN0skddByrPB8CLJ03Cv4SpEvl/Y8fHa8129RFmovVDmhC5cuzeJUWU6YqXviA+h4/++P
wVccgA6YzGQH0nSCC0nZzkcsyWSkXO8HFI5QTAyIfIEsyxy5gmpa8QNlQAYydjymO5XmusNJtajy
3HiZ5kgbIfRmkbEQ9SPiRJgTjO0ZWnmQLUC8DxObLLneXlvO62fRdVLdVjjdjgfSE1iqyD8Ear9M
38hVuBMsKXqCPDlYe+QzPF0bzMmY0Y3JG1YuW4fkVfTZu9VWscf3tIhT8Cx7P1cl7pOGyk+FlSuU
b2gkSEWoapsPfJXTLwStwTbh7UwfMb1IcFmG7jR6WuBa65dySMfRb0f7StFqQGVm6A/iNa6JJw76
Xz3VVaFxhM0E1jz+/4iwvZcKkP9KXOsSBM9Xogu9oT9Hmb4PurVeAOjlek7HRCG0pWYkBGmurUBJ
X9yiTfeEGkC2+CPgyyFzQE4ZH77ylyox2NhZryHUvZ1uzCywemRYLuid2aGGshXy2MhFzzV/VlVm
p3nAs+db1dmWeRRykUxrPz6BCBFUkv7QUnFFqyObObuCCAIqkEr6EvMjE+CEQaOb1esIJaQy1o8I
eVoMj93DW65IVXbChtok+unaO7PtCuqWj8xXSJfLrLvy5AL0p09xsVINmi1Jr+nQoSbilr5JkuXY
OOexQorDPc04XjrX7tqmpHJXS9NYnYjBlTJRoMaZCVT38Vqf5BykK4TxbaYeB+nQC4LEb1u/VuVh
51gYc0YF5p0qbXVkcJjC2+/cGYxYvLmWeK30g9NgKwIAsg99cpAw5Mk0OaK/1Zz/SbBbRVub7nJI
w4Sg4Aj3Cn4gzR2Cxxw3AZ1rPvKsh50GSp9G6MILvhg92wA9KpF0k9Rt8k/Din3xEEDnzzBhuv7b
NUIhGXYEoRXUIDfKj+cMCnNIKK306KwrmjcmrrO0s70CcbW4UElx9ZRMojwJEvZqBsXfRz4lvVV6
WLf8Cvl56riPgdJF+RzIBIqJJCU8Mv3zSWUZzx0ujdyrG4EvjuPmJ+okTe3jiFjBjnBk/2q1rzjm
s74bFbtptH3+oCACnjAFlPjYQYo+VQGMuTbJ18WcHBgR3ieWKYrEQlsTaElgd3903YUiMUXSQgvF
IlShnC98hOfblK08TPLFguOh1bdAw3Kyp6ycBG4mkAA21GPhLhDxFml44zg8AQhQp0sze7wv16r0
DzmqqjHpRkWRh/l9W6xFyhI+pbTVgt4gaJt3Yj4MjbuRmHMKenz/B7JvBuTlcRMZuNmVD1hhZy2H
PuSPxGEX04BbPdZgz33eF7v8dEibw6580uXQP1qXXyU4Y1sn//8aI0NVyln9BQVLf6NINoUbowpr
Ce/Vvm+oabggtHuX9LNMBH4jLaQrWRITvh17v7+3ipE+ybDfJxaGf7cDFmMd+kxEmEMBPYuwvqk4
qa2EIeEWaliDsr3grJJtlTqlnm2uVLNnpmv7/6HR2UqtMYeG/itpY38KQaf9g77UF4hBUasOlSXh
e1DIrpJ3T4qmEIvT6jFwF2Zoxemeq351YRuNscXb385o+DBUqmi1+Xznmm0N6czax9FuNg0ayVYh
5Y0CX4+0KFFvus288VcNPOp/tm0aRJ+pLLK2K2SphCNGSX2tAnzwigggZmcvbF1xUuyHvzBbV62J
iiUriES26LM/rAwfYK+9d7fhNFC+wCrdfAfg0QqWFflPsdxGZnD6HiT4AvI+VX/fhr1aH6vKvkc8
IF6zoTV7JsXJWCFl50RzfBPHpdvGqrtlstg597PsL+Dlp8K+bqUyLJctmnl73yDdzyV5OYAkOpIh
TYlsmtbt85mlkbKuNbkurHtuZ6OxBQoh/+xvJ/vblKrpifBKJpkOgIQ6rjVn/ajI/7spbnQAiVBX
p5S0TMoMZTtA0i/iQbq82BUNRiMRrRzHnLgPcPqDEkUre3bOd+5IFWExywW8XNkfqdsB0+N0kH6l
me4Yrxc0+GNTo94lol7PCnFC1fPxn5pYrAUEMbg1QfsOjBrxuVrJKIJ5zIt9rPtmGteXJXYpUWDp
OFMQbCcFNoewJruPCB5+jdfSGMJ0Xnc2FtGqKhQRVKpwps8H0wedlbNewPlWia3Cb5IkKzPAzPLt
lAXS2eqlST9BGzvRNXUwlxsijCakVgAG+l+oJjlpkNG16i3xctCOlSRXGXREl534EtwLIJh03MWJ
5vDvnHy2WUget+ESLlGclrgKXwVnVY/pHZH3q8ldpqa/LqsR3jA0+SdrGPvk87h16oNPGs5NYEID
MANFd991ty9o0bOXMlf+B7VbXm02yWlMii696xZchs+B/hbNN7KyG62IrMcj6Ss0/E5ulh3Tyx0N
3rQbncTsMJVxMQ4LDu8B0uybWGkvm3x5vwHxM4I7c/o9qhXG2CO2fvOJWgTxoso3KVtaU/fpoazW
f83hpIHTYi45Iz4jDp2zIDgoh5GDv9C8w4z5BOoz1WI6DqbQWqvt2p5yLGD/W+QDYRTIkOx0UuES
8XWPGmG45yx+Mix+1MBEYZkMwPTFxYrtiMHrf8XmZv+viA13Ul5xIHP1+L1PaKlwsHmfvgpBYzZL
hRst+GxHQGT9HzhuqaY5iV0GVO7mbtN2OaxosnkoDvAfTMYQwUyy3ZzK85yZkxnORPEYs0oz2LZu
s1OSFMXjeT6dELTfDLF0F2hwKcW8f2idkQnqR+GdF3pvKERgaJnPrIDXkGo/5apSk3QxJ8KLj8XZ
jteTiSITqBHpGX2apTmWLex59qTWrbb5DXP6i7NvjbPsM8pYPFG6ikBkp1RCeJsBwPj4gukTyQSN
a+R19kZAO3wbKEi+yOLOP7dAvo/RxgJoWcL09LONQgK5D7soH/5JkRa/5J6CcmilcOJL2jiPYMEd
24nE3sUDz28J377LVrR+G2Am7XEGUCEyN2mzDLU78zpZ8jiML+Pmv+OVkET4JotFEIAthoYzJ/5x
iGb5nn8yBv4ZZNoB41gFO/Kg6qNP7JLvtYn9hpD9WSdPh+UyHatI2h4kFw0VHT6zcGkozrqYFYWX
imHac//knfZz6dOmf/ZsLpFp+any/R3JMc32lAv6YIbcgGxCZ86P25IFX24kOmzqY5eBMmhz1lBb
D0ugd3sf6sTSvZ/ZeQt8IFKAeB1SWO3fn2K6q3oZlpDMChtC77o+eq15bu4WWzrSQ84YtBhb5ywF
FnPA5yuak/lfAMehYxEzi87uQ4LF69aYRx/awGpmOw1BERlsvQ7Xp20NWceuwcdDzeepMYuu6yKl
zbCDWSczIN03oFuw78SPelNV+fYB3vcBqK1hp09+akdsutmzhYG82U5/7dtxA0304MTL6YzLqH/Z
9OT6Z8Uz8Td8JEgpgAuK412A1qPbBJNzyUq2KvbJpV4LFQYDvA2lPDmceCP3IUi4fZQTBuSPdBF1
Usv61Ym/4aJL8neYr8M7PV8CdZSKluUW44+qjxPo4f5dpCPhQSsJGfbRs3iubkYa+/ErIdtKKAIW
c5FxQpfdDM72ogYekX0dy6JKtxJvPejwijExJUeZWkPNkIrEkyFcu8zXAbL/+26EbJmSdby0ohby
WqmoV2pY0hJCUjwztnrU4aR/cRNHDDEXm7HlKz/jJ+DGPj7J/rhTs4bE2UlAUUl3Oz5jFHVYK8rw
zYUsw3WAE1tjIrdSrcVmgZJwBjcBgaAgKOX62+ocN8afj8+zI+U12zmH6dTJagEzssM0xkFlTCa6
8JS4QqP5N+f4Bav4qYPge2646GR8E0eQ/EJzxbuc+NHxnXdQG/+P6ziQJfWCSZJOzocUR0SyQW4M
inDLGU7w5Oskuc+drn8aVxX9gf96IWxGyCbl0JEyiLL5w4rtn1eGpmmYvGACwzUv+BfBkZDYvMoP
PyESElTeoL5ojtG+4z0vM9zgfPpLO0e2z9uYtYFcCJdwVmFeuPnwslfBkwMoycnHVaq7Lc1WlKpN
qTg2U5YC/E1gEuV6AKfG4sfdVrdp52QrZIcUyldke/I8n6qXm9MqcmWFI+wvgUOjoktPxpAq+aH8
fbGOXv87nAg0eoYzRax5BE3tLeXAEHgal/yjqx4UQZOsERTDWnXSAXyWrZnlq4ZHyhunaoI/Sb40
s9vqImlwteBlWlWGkGCeWw7X5IWdQY5ULhA2x4vV90tYNQN0VlCI6RyZCWL4MexmyJq9GmHjk1lA
DNVhyHKjtTpxZlEMZXgCVeCwJlUEkhVP6kxYmgHqbHeCDCBCGmzaHyoD7xM7XRwIhnvsp80sNktN
yR/f95ux+WPm7QWvCMtz4WQUym12XX3CH17jYaX+7RIseikbE92dh3UDjgE/8dIuH9jik91phKzh
lSUZXDFhhRCt8a+/819eHhJl1J0IsD4aVGaRdQ28KLSJzEnAHnvtKwLKl8NwPYvARQHxjuOsH7wg
sWxn9TEWNXhO4r2TOqWciAS1eIPl5Cx60Ss261k3lVsCj0DmC24G+HYlm5RJAGmanmWre9I89c8w
9ARBtfU4PDN2jjW6BrvPthYdBPlBSAEHhiI9zDSlYRXmvDR8/Su0/Td/6wZvM4g1rFYGk6d+BSqM
sXnw7ns1QE2ugkqnk8BSgiAWqGbFjjTVBrwtvoyVvq/TRp+GZa2FoQW9Mf++b4AeeagQp7bjkNip
nscc0Lj/y/fpsSbSRbuLbt4+IADXxkNi/gLjE67MaHMoXNtl3da6QyyCfkO3vmrzGaXgRVic8eYD
z7u8FnXhZCRyYX2WfyjZC+3fcxrm6CQ5o48tnhirNW7Zvj56DOblfZ64guL9aj8eOfGysLCzG5GG
NG1n5uTDiOP8CM7DKk9rfsdkMEBHkFsBFf8ik9HPpxSoWFi6+K2mJSXvco7V5NDABNo4RA8XKHLZ
8gXVNUdkPoUsb8n9ESL+r87nq5Egc9RCkcT6gui4ODeN0+UV7QHk6+3PG2B4RXKH7EHoBxRbztdv
DHKotK427ZL29gi251KAcJcrbUBNRH+kfvSkXNx1GVyZKxnmi92N4Y4RtYF8twL5zzWLOj+ud3O4
y13Ys2YBjoiKDBPDo5Y5uDAwkGbkMyl+IfQc4KM3oJDNZElEGXVkjwWmcOWwpt+WbuDXbEYxtuTC
JvUx2ITBolcR5ws3MjV1OmzL4fiwSuSYR+UYZDGnCfnjDfHfiwsgOMOMpNMWDYQ5eQ3vljwbLGgL
bgDCh9UNgKb+2E2oGtmj/89ECViqrrRpqED1rHW9tobXSuNf+iogTfRIBKWBT3zLULK2uvFLTxcl
1qrBCrcfpc/np3aZV1IQuwnCAYV3ZGOnhfRgTf7Hy27sQXahPWnKnmLXj7XHUS2mX4M3wSk8Ayz5
9dHmxPQNxfORHLS6K2T6rQUHY8x4H3LNqv0+kmcUFuBRbkvLrxoXua+GYFz7621/Qt10e+UwnPl9
ac4je2Ktrv2avSrCOJELJf5VgV8XBU1fO9mtm546fA568W76Vdd61Ec7pEitRVdcpVngop/8OKyy
S2mwv8nzRX4krlDlcbZpvZXflvvf6pfIkmLL5wo17npPtOCj3SDbnf+Js8bPsUchVwFf7RWx6sPV
DPJHWxsJH3hFHjmFRLB3VG+q6YjcN5J5+6COjZ1IG3+EralXcBzTdBN1IMYUzhKi+6RiwayDTbCv
al8CRWFfkHFug9vDrQO7sej3PBa4RYwHttPWHmyjclkQ3Lv8oQsgwxAC1ZeQjPPs93irAxYBnXA1
Hm8Urn/6SI4qTsiFVIV4Hb9V6kYMI39tww69R5SAKPBY4NWC8fhKBZ+PZN0/Bsnf/E9AjjRycUxM
gXDSuAF+VsjLaGtk1Q5fnPfILDyy+Jr8T2WG34KfjcMm0d3RJWpggFiyYPJ++JCNxWXqyZF4rU04
6RsOaZkcOrasaZhI6aiMw0yiwQy0chGOg8eIydQjciPXxoBU4jlC3kBoT0bzFSQ4uSm3KFOQZLqU
BFS64Z0o1smXkijyMbpQ+Z64qL2You6bOjf66WdIy12tkrCid755Sp16ejORrcywtYgN00Jqp5XV
Uzxy64RH4VJF+TlolJcMebUKSLq1Vq2mwNSzVVC8D4tw+u51lsMHi+BZTdpT6egbuP1q4MN8PH38
YdK1tyAQtBjH8Z2418nf93qmloWBqbORtms/IAZTjUYkeTYU94mLnPNfB/7HdKREE4WeUKqu0aqi
H49FTf6x+3gkXQUTseugvJ+/a45ZzAbNRS1Q/5Fy9WB2ENfdiqnY66nccyg+8zWn+CZKLtw8l8Fy
hj+ACiAJ/8sxEP3bN+kZ0JQLWLXkPYQlRheO3BAQieWEVawGteV7mL2lfuE+NJR0ZmwhPDpRdskT
Rul7qIRa5C4QihLfbvlwCXpQkZcey+21dL4b/mFJzrw0VIzZDdsA81irICgqVvwpJ/ektwYMsbWw
KJG/v5T8/DJ769w2lHdARSlIKJFt1/6zxrX2wq/zpSVKCCWbS35RUDv96m5gyn9hqtqG46wJNQjn
Unz36dGjaV/qfMrD3Eh+PpHu/8e1Kx2XAatad/NTIO6ksUZnCqsIIVKivvsErL71rkUoGdP6G13n
mGublUv9DcvodPGQPBTk//NFHQJ2+w+hoYhfWkLFojO4n9GXuNNef415LdioR6mzsMqDvF0d/ZZg
1BGbpijcp8Hca+8X0rRvVt55G9UNO7y+ZOq5/7rGfVc2yWORwUAg7s8+QfdD8liDunotmU1ohBWJ
YurLAO6rVNTJxkb6R2ikcWL0hehkjrqROWIiCJhdnyH35spVFOfu/y2B5cD6z6/x0xNawAsPfvwz
SrbNWC1kmN34memh3OY5tflOa/qtX+2+QvWgqfQUeDZnBko5AtN1Pl5CJ5uB0hT6PlbvXrF6JmG+
SPO8Ib7mcsBBKfsZbM5J3qw7aUlMId8ykv2P7WL6Q7fJkvIPAJircea/RQw/9bltQazGusckiX++
bImBYShgzzGHeQHUlleZ5WvkBxfjkApRCJQJio/prd7Pj1povhOGAgGycJ+m7F3pLGkUVicU1jPM
AMmGyI24tRfnzFd1qY7Vg3pXfTNPqGToH2+nA5ECERwm9JUiO8/KCUOVIQRQizkavw6gles1PZjl
a6/aQlfySyqXEDFY02Fe8vaedD25Ad83SMNUh57B4BGT9XJ14oRRlvV8+Sb1Zq/B4aqPGr+P7lzN
0LyhZHlySNTXX23QhYLSWzT+9qEUyjEC5+XALa9O3a3CzEkIH04rzNvjNyRPuYGDLbaCKaJvx4fp
A2jc2qQw4HNO9xPozMyjAxjsw35PoPfgjYKxAAAVNJtl8Q4qqhE7cnmDLKFapyJHulIYnGAa0slf
VpLcsCOEM4saC3RYJuI5xUzTCiaEsWK6jrHmDiI1FgciM/WgQ1L58uB3SG+oeRlaytxnsEXaZoPj
YGBrZl28kP5haRwOmf8cXJAPO+VUvu6iRh4eaCheC23soY9qEUfwNzCdwtm+/XLfuofyQ7kTizEZ
W9MfNfzVxJwNox/4/kWy0Kz4Y4PMx4YlZ96Sux3Y6wqaIrQuHciDpQ+T9kO2+TomRbLuoeClvxzG
WgLRQie30TCMWXQ37txYMeHUV+JZmN2ZRy45XfMEsMaheyRyrOKZyHC5kXCIwuXeSqGwZg9fd3On
zD3mJNbowJu2tIW1723xvPn/rANmVU1bA457sZeBvikXXKE/rXYqCdnpGWaIHGuvyvFvz8ObVd+R
niTearySVq3UmEiXakQIOMX0PoEbuGtiDUqF76E3xdgorbj2IuPf2jbIcUQxc+V1grFK/68YIjf/
DFzb0w8gFfckUZw2Gkjl9BTtnsSigHDPGRiCPDxKxFrNIrOMr4ou915tq6OTzFulhZT60WBBMIPU
OeV9G2VPmk+a6/3QhoAtuR3zZ1QP3UGTj9vCDs1LM6caGSbOhq9TgyVcfiaSRYfR5HhR1Nykh+fL
4xNuiQVEjrawoqPGXd6Azn8U8ovr6NNKTnHRE49FBkJsPyM9yDBtxsOjALbV2JiTXyVkyMC5mk1N
KTKNcWzRK82h8khtHu8CydZXUXmAfETteoxbfXhmDU0q1Evkcp/mqJ0kFekqEdDJ0LI+z0HUb+jf
XCVbNdDeHz5wu8l1nNS3dfJpsAU2+MGo0aEglkwaiwEFv69nezR+K1t9I4ttFzz6HQFt0z+ZIxnI
jDwNRPwV6ZLbB6KCcQf7mKFjJPh1RlfXi1jKMza+zKvLO37KfjP+Z0NGNnhr5Uz11B6YSS7eRKAz
aMR2/kcFKfXp/8qInmTN7EHNKq3HZHLwc4+Ao2fiwUrbaCLSvRPQ+bVuOqQGsYAsSB3ubLmbN5Ep
bO6XtDgHBt83VFvjEyRuEI+q/dESfo0umW4unS/z5w/+vlvDAlenSH7HDfOhkOL2sbDSlW0s3pNa
QpVNdSiLdfaijvG43RiZg2mC11jFTiPSjuf17oQIHuTlU0ZE54Ll7DQjFbO2WG77t2moGpRKWaAs
rMVYG/+vZG2CHFEhcBqxYzR8vxFO9d1lsLwOigwdtj264TOLiOOvvbodyUvmkuQbNI0AACdaDbjk
cV1RGBDLeHL3W1GcWdRTS4udLCYNBNxz23gAsNPgU/kjWk+z2VRO2+1q66zmhumMIx2b9/r7cgQe
w3naTHH5G1Zzja30nUvPTmySG2JTaWMqOXOIxJl0gd+1G42ErklgYAbfZpveV3bV1tYyr6/15V43
Uw3FiUvz4lKH4os5wF9UDe67BZ2ydmQ601lnVXvGuWl+5OHOMXAVplByZSWv0gQ9nNU8k0TVp1/M
G4RATjVsBUOoexwhVvzss4rzfpLkc3S57N2WBFdbYAkPaQe44vTz2kMstBJMLsU6ZFGCJzHWSDiL
TIuSpoPXZhxCj3LrUM/ts2+cNAPCWrDv0ZbCZVhHdzZi1qW28Rtjd6bQpZm+XQT0/bjKJE+iDSFQ
Hvk75197hlCZWLm598reHp2cOaTyodPfFIVLZALr//mKMwYuDNbQPiyUEBkW3YDJzZfmAxxsX8sM
5sMX6pOSIeO+0cBIrEZvg6Wot8C6AlYty571wYlffZ0a1cMFWLOJatYjrxT/pzlNvl561CAEntE5
M+g97bN4UlnhJPPMiMmyLMDrNmpmwCyiAxYaBtDB9t8YJXKq56L0iaZQ+zjwboTqXJWM45+suOps
ogkw6HohGTW+5RsgR0P8bLCB4ASDJsMezjjqoAjZEPA/AqoMnx540TgFFDBZbUiTy5C918ZqyqMT
GQ1mr0J0LMqkrjl3rywZeULXABJSkr+6WAmQ0P54YBU1EdgYKy5rpiU4tgsfhyUYFVirQxnYtCsH
h9llicaXB/kfDycYh58wAnc5Dzki3LS1gquqpKvO+HlIgleCoBzm6zxrNG5zpffww0POEdnO/mwP
R1cEoNGCnwdyAy3WpqmT+oE4oeUJsMGbEf1KvUcETHIEMb7DCo/Q/phMnkX3U+tNcPiMARANHAJw
tOWEwcUpDEakgTtMQNYnsrw0EQiXbJwxdxdlbxmHA6NeeFKdYS1IjTHt2BKWL3RzLoRyFYTglrFD
ZHVb1yCGAvFwZRe/EK13Dtt9qONLljsyCD7AchPZ8pBFnXsAj1VbqBKZkf7ynvWbfbF0V5hO+6EF
TB2WBlXp0yENqaTs7WBF+gEU+Pb4JCKcKeeM5xPCcEszsKMPy2PSPQs+ZN5qma1ICSxfBu8z9vFi
Pyp+auOoLTkt0rBkEK94h/k0YzzXAz8eZbchaNqniCTiFul5Z22OEaW0m4FC+jJBX6ynJCpK+Y6j
qE+UhWJTvs8HCChQKur1yhsBeh/fYPCxFXFvAWaqNvz088r7FJwgRx3rEw+X38dNbQglOXd3QM6b
hZJlXfA7++RxWqhSCob9QWmoFr21+ukJANEzf12B1C+AtWGsoiTwQF3ocyBbXlgD6AG55QPX+xjp
jTtFP+jY/zAUIhBbzBDFMFfKjY+l4oE2txYJJhpHne7av6VuVdu/6NZVgH+d/6Z6wVeyTC1XO3OW
ZAQEZwTrF+dfCF2lprKEUg4ZT1z272m8nekXbQUK1cXAvLfdK5Lw1WR4rtD6d7ctwmKmCQVMv9e1
wf34DcQrtu3aHIPYYjowAQgssRxLcGMCUV120y84vM2VjOHrXAnksxzqvmaug+q//pTIS0xZ9Q2F
VbaGYDN/oEId0netPADN1479b7r91AfCs61hLKHuGqN2gWQLC3wVIrrVsQKasO0eHL0YJQfSbkrO
MEBEWXUJfrlmH4nPUx4k2U/xz+Wi3TSCfgQ2G5fWOjonYekVFM8W2tv1ewUEdCCVhS1oiXnjnuS6
uEYuEM/qjE7YRKtv/jGBAWUFwrGBldjfnzq40jy+KsKXzB0Q+e/DS+ZVqLAfz+bIpWT/uBAJrzS9
7eAtlMDOqeLsyQ7+sfxDSSYe//1ywgyWlsNxEV58Mpoj8iLLIOC2hpwNXD9DdynJpXDXPsYnaKoH
S+TXsyMB00xqKQ3O4RQ7Vpvqs/wiePodETHe9zFqf9gblL3UcS4FEO/lpVWBgiNiv4wuoorQot2o
hIqMVrbFqVBgdEjhyzohqTrhUlJ2VTZaPKYy6lYwRC15JRShYNXMT/9fibTg+b9QanM7D20hHGeJ
vUW3uImTCsKOSHMgfnGBPCRtxhXDWKs0Djn6ao7bTuJgWK5KK/VF71TUW/wxuNTfPsQPhUuGocfS
eGoO2E8deUnsHvt2ihCWnE7CW7LijkD310L3FqASZo1j62XcOMDWfcyMrHN3HRC8iqfg8DNKqfwb
px0muwDJjbOJl2l1POZOHWxVFiyhmQNZaR6xWapAiGIUb3R0muJa5T/PU5PTQ9iLnZJA++3nIw2x
/uJuLvsL68/djMQUb5XXmKwMpzVN/t1PlbClIpYX5WTyKAKNeun+FoNs2oTFh1JMYGpeUB/mR+HG
XUt5qUAqYiOGO0Qdy5jV1xIg98ipvZKtvK/yARKZ/vKBv0JhcoAIazwo9RYJAZ4UwoqkBzk5nfsT
tbmX/Sc6VMziBWagU+P5NHCaVBvxa9y/JhXVyMfHLQuH9yJV1Z3k4GcS6tFgw6roBNiKAXTobkKW
x8SIPB5o1Sz6fyT4GqTu551XP6O3gb91HMjWRA1rlk9HgaQrjEw+0dPTkqrLXZrxOtf/kFc3Y7iR
MDTsBGJ5heUXsJXboKZYC3c/1KNCqOhp4XAIYoPRP85iLld2ayRjsDLIVxw3ym/lyQL27f5NRpIk
XF6MJ0KnQSr5dOirdkm5wM5R71W4rvP5WKVpFRaDqeygo6RQ6Nm5Egcj0AzjKQvHvHs0WMydXHpi
29xIW6v/8huS8ZwJWLCdIZrkNRSf/w15/iz7cel4N9KYRelKel5VuPBMPGYq0gCgkO9+r374xhhx
QtJ8IEPr2MrPs+w3ipqyKFP0V5tzPhn9vsskf1ZRSDqsvD+2nhPveMVQ+7bpGkLUHs7iPIsWuWWj
HDCuDv/6EwstrXXGTOcg24myXFPuS7Vz282xqpO1soj0U9HQhFSm/WV2y2gMjwjdzsN1LxY+Dkxo
W0gPOfVFgaKDlheFT19EOZTM2OJuRX3geQbvTPPZx4QTGjX7Q/K0NJ6MEw6MZ8rPxuwR8M/hZacr
RRHrNHkMfjW7ZFlEUplkFxKyLPf/tQ94Za3p5wXVnqz42YfnaS6wRyuuwtDZD4llgloJRP3QO8ig
xmXCuGHzjykQa/FS7pPHkM2Xi+POOgPzOdVH3CLZrLv3eybtnBZPf6H1vKyAyuQDv7vDaSqSbiOr
YXUxJN+vUUjCdwiC5il0JyTxsGupKW6cpXuNbeBclZKhyBaXQu3neQV5ROHCu3/689+KZ2IiZeG3
EpP2VQ0nzaat/QfVkhUbtvqHIG9wZz2z3RjGKnTYIS0LX3lZGgBokAJFgxKZZEFWHPMSC2JlKScq
4r/LZ+uuhwDevUK4C84jJUVA9W2aheFlfwgWYUA8Pf5VPVR7Ljtlp3nKpoMqJsgl2eIUhLQL4Zjy
JO517izPVuH1HW3qrCOiKR85WoIxMOTgRJ8vd/0ne78jVLnc0ibDsIhBfQzrg2FvLFhTvSbaFBTh
4qsEh9PJA3L7Gbd51qrJIyt2iZCNToNUkG07sgsVs5Ojs/tQqaDBAUshF4GAHk1TOBrPpXkpAGf4
pxAuRZCnR8oZWNzf8E1vTFzUF7yzE1Vgs1HWmGPTgPGEexmUg4KWyvCMiYnwBJLc/spzqPsfoihc
QWUSYVmf7FenJll6eHpkJm6mhrXEjbNlb7XkXvYBbB5rCFy4DtECytqmEwc8pHe1tE3fEoZJ81gF
YQC2JAheiVp2LeOiKpThKH4VdfbXl+WjY/aWYfrh+yWa9YME2Ey7QEJFfIMBUZeoNoDj9plCga2+
yuXU4yt9UqwrQ69IObjzt2ONEogx1Y7wzReVmuzLuE8eub3jIDHGxLJLeWveM05Ybn1nHE0NThuY
9JYEpaecxOjchxgyEBxW738skHl0KcNX+uMgkRLxitG++TsAdZ9x0j8ty8L44BxJ+0ksMrKxDcUA
rXVR/u9aEesb70hxZEtt0FxQ2g6mvgG1gdyX4V1EzqKFiJLhD+3ugOH55hm8j8MtkuHfQTTe9qQk
aBQJpI5lJDT3ziKBjEminA7KwwY4sKh4ffd8tHWZJ5r3wBcD56EOFdkxSOnikiBTzWgcHdwIjxUG
/98L7Xem4gykyWLL3qJ6ar3XUB+CFzEyPeXtr9h3LoX9v6IrLd9LKoEgA7frjY/N5fdPwb60+Qxh
ev9YFUHstIdVsZ3NJGVfJv26gqUSYvbRYlGFZaoMTuLK9MtRr+3YAerhemQTA8bpDAvi3dsXv9HK
f13iD/W1lKROuLLKkkp0rydV4e9FK5FXT3PsyMeMrlW1XJNKOyozc3VHRy7ecQ2uX+kbqUO26npx
XRERradpKA3Dj1cBmeaWROdeDNHuGx2sAVtFIuyQOfkXgPIDiDI3NLcsYttzy/dllCkUAMSXTrkc
h8uEoH0LeL1BbZlAzRoiGLDNahDlxaPu9CetfkPR5HSi5QlldjqqriyokyiFLQZ3eS9EUuITyVcd
mofmnMf4/Uu9aMbIF9S2rHPImrQwOVsYWcIeeVbwPnKHVmb6LrNnLDXuE5zFnoKiVSgnk1SHBZOn
YyiFa4pPzfDm8SAgDtIgYR8oR2vYErObB1eYcL6VeBSXq6ItiKBMUB5jwmpqQoWxezsnTEfZOalT
kyuZuEkItrqfgx6RsM/a0y0jDhgjPbIBdHvXmk5ejmqLv0laDWP3QXAz0NUxN1J4lJ6TruPpHIdU
Qv0JRf3MpUXkQQkRJuUzz/fCLdqcrscSoCvuvCv7cQtCzo+FHJ3IbQCk96bkkP/yQSMR29B+3c7q
BeJ3GVBz3hgSTCBtuN2DGyqCxRw08d9ANzttIh13QnHel0dLsZ3ufUAPvOK/C7kviZXXcpYW3TZ6
OOxy5jhmvtibuHT3KD3YeIFot41zh1EplrCVL32UxdBkUu3EBTjE9rLLcldlQVI++rF6pMj2xZvv
IDxsFFft6pjbMDaKebPWp/rRsOrHm34wB5044ENJpuikPsYKlDJq6S9JTOzq+qauCCXUcY/4vTQS
zLGa0GxPoIHUJnV/5kuseTiYE8Bcp4u8nRFW6b3xBwvFLuecHhN7Bel62hai/6AaZyZUF+cIgMaz
BJ1+Jrtt1UntkcnfuYfXeZon9QjVCoFaHsciBXm7dEBtE1mL9+kUPY535ZK2aB3wTFTvnSnzHyvE
XW3YocFvDIQsyIOaRrwQEdmmsHRazQCsUtwKcQ3SwLTOdNG3SIjgbNt9E/U8kMNJbPeG8ohxxpeL
nxu7qrTvgbZis61Kg2m8MdbhxrXtTqsEw/MbbdxUWhDTf2leh0zNspp6VHsr9EKSoei7jILp603G
/A39aHFORb7Xd1m89ZJWiUl2XPXhkm//3R9/y7Q+jqAO3avSS6t2D5KOu4lh4XJQtLo01tJXZYj0
cL+9gyCG5VUMuiEAw0PlRSyz7O+2tMN79RSZKrQqd3/VMiU2ei05NzAFTXhYc+F2nT71ChlrGOJr
KCO4nqdhrFlR8rFgfFs0UW0UQr3z8P2gR7kgWa0Jrmu+72OqqiF+blwLcrO/ZkzAA+ZdFVINXad7
8qK7TKKtnF2XornKZz7XUhxn5ztw6plGV2aeG6+9Z3Y+iwRjccOnjT84dVLstJleaM6Qoc17RzBr
Thy3X72xkuy3eNPz4/I4L/XkhkDZwADHjVlIQof3NqkhAeB/Gi8Sc68jrfjxHd5xpyc0YmPhG+gU
TKhxjTI+24A5D7ZUf2pxAR2VZiWDpOaqyItr9+fnSx3uInz0MCC+mt05KaUg4glpy6yDrBjGcIcs
s+SRlHJaPyLMa/m0xuIr1SUGe+J85WPNQD/VaehOeiHUSa8M9QWQkkH0jhAeI5ZRtOB9FcrdZK3N
4ygvv7i7OeOCilRYJkz3RCChexTfyIK36ig3rDC5okHNbGSdBKbg2Uikc3Qzq7qteuyg/HuauVtK
21/Xq8NrZtjrK4cAIN7CZfSMvgerP57LDftSPPkrBZeCmFxvgczrzG+BTGtNXazPHFVBy2KRuN3f
btlR0zDETyqSMZLPsZY9Kdv/k66Fpsug7Q4DzQhYxRgWwWEz+70QR5+HB2uQrfR4IsS4Jlil+kT6
NAu3tiRzjZpFVfqGlbCj3Q86v0GEaI+TM7Udk4MwpnIHsvWYJmleK/F2hz9AOiox3Hd4RsYB9E0r
1eEse0o39dCb2HSq0S34QEeFGlZuUZbkXencuB+Is4I9oWHb5uQYUVa/duL1exG3kA4E/LaRiWM4
aYGGrSUQgNB8v6IW/nZpxh5JqC+wxvs8fJvMQE8JpocUTd8nwxIvAg9NJ4lFue+1NVNaIWC5ijao
CH61D+p7jGUemJVyyVG7zYPzVViqThtDPQpvh26TYloA4Xf9dh286mCvER72AFvHRav11ChcZMw7
+Iw9Hm4vkXxq+8bFNEpGeiQwjhx/MNjGzVy5QdQJpAoj3zCuiAN4+QsFLAj9TXS8xYmIh3FCFWxt
F85uHp+x6z6I2MTBXkgRfZfOLUn0dC3JYICa11HcDD4JKQ2ptpWjTn9oBKpII23sVaRaKcOTpv1r
CVehMj8fgoYJ3IsaQY28+KlPyetp7T6E357y2+n9B76uHr5qElq3b44YLiqQSjwmfRY1CyHCk+4n
BIuFgxAtHLNltlooQYfRDIUCrIohNP8NxDUC/6SQqVy0cMBNq1K3lh1E9zppuBv/kzj2Ie0dWHxO
ON9YAJSRuTxP06MB/buBleWQiavDhgDmAiTTin50V9TJeU7mxFkXbx8dpM24Rhd16h32mSl9fmMq
LXkAR7X5wm523pVbYT9IeAmAmZUf99hmInlLadBX/6YG1HTJbgPBo3tNxDX5wQVvRXdB8uUKrrzw
scibAthSBRePKgiD8ZKXWYbLD5gvVHgPrwSGQAvsQI5+zE6Gxq1ZGrAiNZ3cgcAU6wMtIpCes0zy
0n4Ewp+QREqa+bmKxbRLvFZUXukqSn9sljpEyhhyfvA4zT1xWslQhLEAOcgRhIdjZFfljKaPRtwc
XH2QTqIbk8ekqTvgHIkJe/TlnpWDbACzFwwEzxfZTPAgtdycUNqW1Ya2bvsrSMQ3TEpxwYIP9j7o
BEMOqp8hfXph68mdmX7kJvX1MmW/vLubhqwvRjzyAfsqdHTczl5EyVwedzl1bjbg7rNgvxcFZyLw
e2xhw9wq6BHfvsU9L6cr9WJjNc1ZOiZqRs5hwfyHQvlmusKT4sbrA7aHyIvC3Gme4m89I5o96cA8
FXMGPQY1MJjqjPSuByHAaCXt5yQsBfMoY+FujU+zBNxhiZcWoS2kYo0x5DpC7Am4XyJ3IPYyWZgs
ECYOfcH//yiyZvUTJIgpWGGGuDxmMoekQsyThwaR4thdZsKUuADp6g56l1gOs5GUMCbZfMs0skbx
KjcnjB2SNyq5m5vlEurbDRHAKOYng+tVLkrijAWnzMLdUlXDIo00VcZfs506ojctzIxnKez8tuce
oO9dt+h3aiiYzvSE7IYPqWX9eC11khTDRtZOqiSj9EYLzKqi0UI3OCsaGRtWa4Hvz+jbtpPGU1Oc
i+npOZz3IsfDzOq7oPfIRWYfUlqzALxYsM8b+PpJjecsjOn/sAH9H+sx6dXK9Fl+QGDTYM+ae3rT
zCgH3SoqsDMg8U5FG7Ydfq7ZgXIIKLT/bOHVjMwVZqTlK9LwZpscNJQC6uSDMPJLJ5bbPDY4omcN
LdCVnF+eZW2QejxUwol7/9r0dO7jeDQlbEsVmRRkXQC0FZfh/I7HCP33XulWexg4qPiF7punlGkS
OVRXwdei/usPV28S3nEUVNKkXUTFMm2CH9tsprr2UblhiapEheIuFC9u5VGxcu0m21c2D2AU+iQj
vcBqUD1T5j6Q96YkQy+1G6kO4joeWw5MVxD/C+kYF0ttXvQthSrs+0StdXlSPOutx92VZ2+eKLsV
Dvhbhi2VGKBvBiAOnPEaSDHot5wPjEObnnxcVEJSMs2ccfAZcJt2cFBPK6xr7AN4cfop8VI+/7sM
eRgtLKsLl0ARCDrMlV76+7cj+FepUN7YR/470dxwyyHdyB7FNKaIdRhLsbFuzZ5NazR+XinUyrx1
JTWqtziC5tgmcylFtCyBgovezelrExzNusjRjSFqk79EOhlr95J3lZFkyyD/rONAxdveKDoffiI1
yyApvbHZfsgHkO7jIWWNgI2uwRpPxtYIY9/2/qYnbLAB89fOuEv0w4CAh0SuqoIVRV9UBY2SFrEu
DroR0CRPliz+VzwlP038rfBhABrzv5wtASqjWkCB6E400t5ZgNWITwS1oJKhgTqxG0LhMs3cqCug
3hHVWn+6uwxYCEwTSssGSWRduYDNf2mfHmhb+1uc0VOfXMjm/RUSaqrpIHtNkaHhTf3GL8RAj++R
1f5iSFcYBTLjLfl4IpMrp5QY8ezGxvH7/M9NAyJ+GcyTs6TFT/ANlibcU/W7b9G4vWr6wQHyYbL1
LKw05i+vxQX4VVjwu/ssccg12eh4T+HNm0HaFVx7v9bMVPR73Y0F3KZ8zywDgM39xb19v7suYngZ
DqD3Vwkn0Zkf5oEiptGcGHLBhuzSkmaAEiYDMl9Qo/TZ2mmBDl09rafG+ulpyFVn80pkUfcF+DlU
RIDyarjpvxPsM8EKkcljg4/4Jdza1vTbX3JW9U3CMFRK2Te0M+OanhZWCI2LLJ4VGVVt8DtcGBbY
VJZmup9LgRc7Vdos4xy0FEwzR/1Cjog4BXXCWnv8KNcYKDyJ2x0q1zAS5/WAP3QiqP1AxxxazMOe
3Cna7u8cr7IKtb2qV0Lg7tx7Mh68TSFv1BCP5Ho15W28pZuggctS0D7/bh4zZLHJCnqnvr4juRzI
+84Zd/aHG2IHJ4bhC98HpPKcPLTEbvKl56QoSARWVyAhQvDoaYHdcuKOiglA+7DSrMki8YmzfIj8
s9eZg/Ntc0oF/VwHvlQLZI9oBh86YFYVdCLmkPbob2I+lAo4A1bNwdvISIjojiib1+RT3r1Z/iFQ
lmNAC2kkni/dP3Z9q1xsuxmcmp251lUROqWWx+GFrY+Q3/cDQajXb3mEEvTVpj1Kyx7h+dDE9VqZ
4UKkFiJWpTfxadudZkJliswkfG4+oRTDrByvL0UCxYZCsLIRIlyTLOx4w3UdNXcVRgSErJoPS2vv
DM4I6tpNxS6wid6nZuGom+DSnAetsmR5qZosMi9JqLH/9H+3gNj30Y747UdRC8X2GdarjsosANrD
bVbtAhKNMJ20eL8VRD5SnUqTVSC4AYH1z252wVmEHJvNhlUjB/uQWNgR91u0KzN3GmU/YvFH19w2
CTgNGZ5v4MqIxq/dxGMWPO3Ty3zIkiuLsHSvm8ZEDL9D6u6FvC8cK3jksi/G5wu49nocArg32GrH
bK8T3zTn6idoIwDKRj+EzGjUtq+YQgDP46KH9e4XxKZK6a9Gw8bpJekApmW4ebEjSc/TKTGaQGlS
clwGDh4cpy/TgXHwLQvLZ4i7pYy3HIBMUIHlV3iPqEhwaU2Fq8ARWc/Et9DfW9N5UzhAK/UZNOLF
5YzYfDBGN0KnQB2wwJQdfV+NuqoVoiYhEafLVsQyB9PALU5OxekNfodOSnxoW55XJ38HM64JP+rJ
+p+kNZNdBLuvDApqWzKM2i3SLcVDiDWhUH/icjq2STcdT+VYhU7Bnxr5DGxxnTAu7lWRYYhtJstN
02Pxpc/rf75adT1l46TIPLbvm8JyMAZLUNljOcM2f0wZWJApRpWQOWqMbt1cjp6+hRNOp99veMGV
LIrfQCtCpHY7CvikmU01U7j+PnKdzMNVp41ebjbb/ky3lwujTxjjq22F+t83i+hZ4/aIN4899ZqS
I2S7XoDyjc4/S7OXKMGa5J6+1ITACWvJbakpN8L3nEosNT7U/Ly+mIc+ipFaRkCqEHpX5d/w5NmO
UihtsY60FAlOlCU2CY/GlwjDpmv/674rdRRKSSXIBHb7N10+aRBTv1HzgqTzsrcsxwqF4QD/8rv/
GywI14kTCfLJsfNsx4JRtT2sGfP66oC+/y8J/luq8vmFH9/fp3ia31SWArnJAnay2UEdNHcfOG2b
BBvulox9lLqs1LjReHsbh5lWvfF0jL4FejURikcmep2PZTruPhefLV0YguNAU4u2yanGRTGvRnhf
SRxwOK+OPNqJeXLGV8HL4UvDZdxzuWRPdPaWSyIrwoqAP+nCbQ6Rc0j6v1nIWM70c/chDDcje4nr
g48hu23ik0QszSJejyUqV1dDUs3Qnw0+ob2nVogVUI16/32JMc6sdk2Lscjq+FrrOUMJgkX33WB0
ybu4oSSifqscmjpUyHT+O6zMe1FH0l7myJWahV/JVDgNAQcgDGIT7CyGnqVYkTXfRPffMfPPOgs1
VpYopVPPYTOy7Txo9XNgzB8ZtA6NWhbRL/gpHZGTNwVM0iMiNbuWA5JTV9GLFttKHkFoSo9EG8f3
rf1zE/rP9IiqSjOK6levGlNGWeIH1NQCD4yWkSKo4MZ0KmqhqFSC2OFuDOlJI3ac4McFQaMzsyZU
PvcJqa87rPHxB4nAAQ43xFiLpwpzZD9BS6b7cxIf83FV2KOgCsc2di7XdPpRnKqOsojrRzcNZfsB
3S+dWG/W39kTBjb103JSDbp0tXq6atWxW6dzBzWhmJb/Vbikmo4H8edlBWlqa0I9jmzIRHJkowda
f1+lZCPlmwt956LfqQyMovwTfL6zgH80tY4sf8QGaJe3LV9bsUI0XcW1BsQos6wsk70JAZK+6xy/
5Ma58Mqe+JkDLLAkRhGwPAgS/3u2hAkffJfgkG20iRoRk0BnXO5rU7SIPRdkLK9LzmubDa9oZLvr
Uh1p0UIvVvLLTx1+EgmV3wwjOfRiKLLo0Z1ARIS140IUir5OanCEIWWZKRBeAff1f8SkA+b60Qi+
UY3r50Ev8EQrnAFvFeKzcaBxdMlbWsoyL7BB9uHmaFgfYguF2DLumn/keL6rvIUJvlZlLA26cjCI
xbDq8VQvo+LO0nYa1jt+rtIpzk63Cj/D8Ky40oczt9xu3qUnoztLKRXvcU157B27AISAlT/n8zPP
kyAr0ug6dPTLajYiRgp+xh3S65WPRFu/MlfPf7TiALMPcXg8Ji3ZZBqwIw2QzKzi6/NzQAsB4g3O
ixxwMunm7mygNRxCI9fLpvkOxujX99skAOmXYiwnxoCbvbdONMfMn4QFvyjF9qMmx/f3TAyPFuMz
nWMZzr2iIq6tlYTN/i9XOAPPluEehv3KYdTQKDjhlYe13q2faBSTwGg0vQGTB6wUq5fLkcBRZX3b
fKkqDOUpjkkJ7bWx77O2hjJZNsuvNPBATK0h5mdq4MhwKm5ffuDzWQPLasZHP4ISvbz3ydYocJSc
8ybuVKwkpPgBEh2WAyFRBPbs9DUXwKSiFgnVYoQw1z7bBreljeDNSkM7AXe/o3ciiRj+bvTcx/7i
VjOTj6kPtQ7yKnUqmWg5lodMqMzdkkt94KXRbHmqIE4olbyj+FouXzRATZFtn/msaae0odD5BzEC
CrT7WDFkLdCim9HbBrCJk8XWqExS0gdbw3AEcd9BJKzwbsoWe0vcR0Upyy7eYiLdgKMtkWZxwqpy
TYnDeBE59pIYc8lDkA/9lTjJwtPintOdYAkSVPB2hFEco7u2LzZpX3vTdBGdBRzf37Udcbn7nDeJ
DLHGF96aQvd9lTSiU8qQ9WV/yoW6aIgMDX/KdV2QTz7MhKguoSSl0REM+iroA2LYNCzpW1VSWgsD
hwEHz8EMDSbuZyQA2ngi1JKhvkYCofyNc/fRkfVbk+cwJ7CRWlD/tPWzDMn+rTHbzZVmZdKrEylA
YPIM6Gs3LDV0wx4GkAmM2T9UpYufGEjmdxnoGJX0I/TdCSnE81tr7Jak7XbWksAMy5PaITRYn1F7
GSzxzq6w8GzkN3mcHN88CatB4etfUJ/CecN6U6EFNWThw9xOJPofByiJkjkPoVc24iFDKkALMw/j
Q7in3G+jEy6LljWW8RAFPHXitFjoM1FGPGlTj18/KEuisV6TJBwFC3a3Ff5MMkBB1UFNwG9B8OQ0
bY3n5s8+M4WYi01MsLj4bcYNvsefTx1neEtPNjtC/PnxfYV4IOnbZ6HU/3D4iwN5mcBQ5XnPac7s
WxwSywSSVj0/cyweBRzh8AKEaS4fTh6PemVjadmY9NXiMeBhdOik8QzMwyzHUb7/KHQkWWz5h5YW
osCnASXTn8Avo1P+SVCK/2EaJrKWeAgWlHdkG/Dg74dWbo8DlNw7CxpMM6rizyyQRcKzg/CX0uzv
i4cVlKw6QjSkWIOq6/K/MxSlDx87O6mlpNL0uoqI7w5B+h94eTxMqQH66b9YQ12l7fecQmMUML3Y
qQrfqZJSZ4ZYzAY1QlM7KANOWjAIiNSDUS9IefUZw4J0UQMOCHx75awR2mEi7GdzNGoDH7dsvXzD
Gi9o913SCkgEcA8rly18L5DFt+6jQtaFTryc6XgA1KCWw31374mHrQxTpJfrKC7EsJ4CSfvEEc5I
lHHFwoGBDV2mjV5Zh4G3KJqrQeHmPCZFJwDD2uXqjdLtTNu3NprFglslEGtlB9cFse39SsCj0b83
78boIDgSSIhQHOyLOvlc3pY4kBgEYmPeGmmjMFUuTj38TwDnQPWObj4uowaqLUKfat2OXdmSTDcJ
SeOXbTKA4cwxuyzzQBOBntcmewJznchIvmiZcMa78Mz8qM+9UC3F/0qWMuCT8im8uPaLBvkqqvPv
16YsAYZ1taQdG44l0MHi9OVZly5F46kokmOCK/aqAwIMZUPiJ4PeWDiii7iZBqFcX8evsEWGXWmp
htnw5rkzl9EdlvPqh2d50HYEzUmTsGJkHPyuCe05q/5ffaFYSvoY7FxxTj8mKiiaKDneq/voIYFw
x3eU9Iqx2geUsntB7VkTDG/qQA1QSIlBwQV/3PaCH4gKny96zYQwbbklN80m+TxCsliCVw7S2Mgw
ZN7UPJMelEIyUltsa6psrWXUyMDiHFIsiGKN2daxhEbKNhkH6PZakXW4cT77GOJql6IcwenWvrQT
5lh6YBJWxQalgc1rjmYuG9/aIH2tT/A9OiqLQGzhtlvKUZeU3nxm/sL8fSqmoraqbT1GikVzNPQq
PoTGtOZfvzfouV7wOEPQSA7fyceH6es4Un/PCF51vmryjW0xnX2lhYLny5ZnDyroUUN2Rosr+bo/
s9g5yfw7cybOM0+COwYD7xxkYg44ZMPy0W2+UasSJLYOpcVCkJMO+ejClx5LRoy9GPeUDSnqXyry
pZQ/lIFBLxQBuj9R+QXHkOyIU8Fk/76UM6XTr00zo9vrn5yEvjzCvbR6ISlgXjPGlsqTg1UHkbKR
bc6+hPM+BYBI2iTHxq3d5BSPiWeLcpqClAyA3IQOUnOzGgaQBKUoPAA67NGX8eqF17Q6uvXlcmDo
TpqE3tc+hph02ItzyNlbtTrl9Q6b33F9dZnclyh/x30XN9alP1+XRv5yrb0Hihzg6rXJ/TKS8vtG
UlUPgAfnEE1IAsGnJ99lZDGEqiYay/2xir0i6H+BpHBGoNzQnioKMLTmaAJTv/W4zcmd60eDsLqE
+/jqgVvrsCisPZkId6gOgxIkz0ooOD9VxwVS/SMd5rekQt5AWNm3qLQgH2ezdCSwVm8dg66y32ik
VL5w7QJpNfMvYOW82AhkxnKIYHXWI65hCaYQ4uhiURPzHuCcnQLBJjzyaoslknvLRF2b32Aswky7
0NVVCWCoEUHWjPXpTa4jD8pLdV36cXuduGyKvaIeXbDjb1Ob8x4vLEoJlt0yUT5UiLnJNTp0A817
Kn6d1LJV5W46p/l+OD7hAKX9frYMXVBma7l3LOtY2h3VVpRpGOMMgQsWn0uUmkmMSxfwHdsY9izP
H+Ykjtx/crL8WQTNIvQIvoTO5IRICn2o956ALQaXzDaUELMQT/2tdt6B199y+G95VVAkXUUmrq9+
RBUc4h68IAl7Dqk/ecYbWVo8iPV7Gk+NNU6WaycISwfHnW6hoVECux8tmbcgZ6LLfy2wnmyYUE5W
eF8GfI4lHayJN7k7zaEmkFPPCObVeBMiJj//whlAwwPFcDV35o4TOXfXOzkFapCVpnqV37GFufCn
lncg64bDKdAqbnjDGZmILDM2peKBoVbnuvUDK4nHSwe3W0p+bpkhnqJZYLs5G2DAi5U/827+68qQ
/fdo8nAzYYvyVqRrCxWar9fdNK76xisyTPmrTAYv3oNu4fiRx+9i9viTo5+aAd/07NpiYsZ3pIoD
0nZPE12x/nG2nr0axPcylWFm7wSIw+CkKQwft2neL01VPSi8m1OgKY7hbsToVmwJPC3Fz920kkuP
R7vX8KTx6PxnB+o5sSHFDBd19scLK5/TH/ir8b9cpuurB6sbUD4u1lPP8cV741hl5GgYnlAZWi3S
OpAWDUR78RZiVypvaUplLyD49xu5IDHPwwDrJvAj+bd8J2H//L+Ss2doq25uco9bGXRRJLEX5g2y
QUeGUy6m4OwJ8drlUY6EiuSmVA2EJdPRtkeyut7mU6CP86ZaHYqdJCWrVKsMVaZBdJRF0xXjJuCJ
964KQQXVtRms3HhVxmsg30zy59/7yXOqe0GncYMFH09HrgXfe0IlJvQEEp7+8TPh6TsmpDBa+2pv
V3501byzkS4KNZiDgSKm7BdXvm46z/7q0Mn0pDPXzZUl75zZJoh6BOVEvMiupqSAa3QdhYeQJk7r
iLjbtTBhirSBjBEPg3xzsLSLAdGFB9Z4Md3DicZX+u8lwfZpPcUiI2EUHT3D8RKaY9NUhD8I3Vr/
0U3vIknjFfSo2TDwjWt13OW1xc7cUW8JorZjO5zTV+cf01NxQwW+rJYcA7zWzb0uwRzrQS/wN3gp
VmJVSt4pkDIufN+bKOWn2OBPc/iDGqf6ELccgSzwZtWx7Yb1MiT8lYEpc2lAxVtAI9Cc40SGv1rz
IjYpNwxFE5V6v+5y/oUSoZihhQEiS/hR7OVNVmoLEFCXUVJYrtAnkpIn/+2GlAPIssSJWMivQ1eH
TC27LRVFD2kr0HQHD596gfkbMbYG9A3/pqKwzHJ7qz9uuoWaJltP5L9zAfwGX+sMJTpJ/GheCEFT
MDu5ugcF5RkIyh8GF8Dc2kGaWOI26IeYWKsmNfKUdnKjGoDchvwT1wAgSs/IO73LpGbj4rSM7UvQ
cq+Hn7vMFSfibd2di0In2tL08jRP3nUkwE3LWPiumH/e2dSuiNq7RegbdQr5M5s3/Jbm4wC1EIp6
BrmnD2M+ijtIcwLdAC64Brbg9ncVaSKofh1XNKFnyT/M4phlHaoJk8rHw871BLjuwbeZouPrFwth
Dsz8XAJ4Y/QISU+D0zc9rsHJ57YAiJn1eEdlLxhIiJoYuCy4DP0wzK60f0ip2C33TA+Cwmta/p69
yQea2vCerIJ2Hff9xUvnzSZhl1jmBYw7QTiOHC3ZOncGpDIwHROtctbOiUKJhyydTacoQBzFq7JG
UXtk+Bk7Z3Sx7ujL3wqMbEFm9Kb5sPtjocObWqwfWr7uLEevXmP7VKDYnMl9cVwbeCmMwIzBOsoK
PpKYGlGjDZY9N2jM/o+Tmj4Cq3Mbfam9tk6H3Fm4LR8RiJin5pjRnT3RQMEAZjlSq9HBfYrca322
ep/ijrJClJnZI80YYFZU4hSonQktd/qFmd2jZ2lZVNabpAOpKPMc0ZZv37QNCHYcNddIdEx9w4qf
YwqzoRDNzRY5T4NlbH6o+rpP+1oKyJBFdLe0zMJD73zjSe8yKOHbe98jt6dRvnzZxoVP6L8XnVdx
Sa1o/rBc4LsaIFdcBBF+2eFfGE7y6pMLyMMOxbgQjAOgl0YGTjgt5ZTlilHBtsNOiO9wKMSb7W3j
FEH398ebY/ova2PVd6X3n+qMX9S4pRMqdhK6SpghKd1Di5fOvLZRqQ7EV7eoV+qWfu1RrP84By+Z
7BUv7f5QBfgOGClVNmhwpWUQVTp0Wh7LhvVwgciPVA4uLjKspuCKrIOZ4GIvUtdzJmGWN3cUezPc
jehg+b7DmMf/WZJekhsMNGkekbLw+RyQZdAfnzXCLVmD+bTdCcVi7c+MmRbmS6tSuigFxquyb+rP
v6QWnLbLygWlLFRw1Fa2sbk2XNKG8iURntTZrd2UCQsx3eVJQOBNfhdho46uSdgVXLOIAW9O7pIL
8+0XqbVzXtUBZ9nKgFE6s2ZJGWsN1dGMqevrY/ESiFmGodZwHlxrKWN7XrTlnR03U1R6nlo4ACe1
TvCMhy4IHhpnbcwBROYzTqiHGH0FjdfIYQprJIIefCCGaTl0GzDVB0pzOdHiueHR3Pz4aaMsYK4O
1y400SOtb4xBsAUAOUftMjswd4IMhM0fTBUi95tCYAqqyo8MIvAdP+rx0igHSCKccedeRZ75a6p1
f4/wIJJRLXmcebb0mJ0J5YJ/fWSYvmmjhdjsWJ+D0TF4NE1G7yiMopzR3hJokOAVYdV+0c8Q0kUb
napaPOObZ3Y99XmG4Nr2jJldFYgIfd8ZVqD5t9tcQ+t04Qbd/UBf3gqNlZ3AU3CbNugxClu1BYNv
qJfP4BwkI2HJzFl5UjOw6flpD8oSmdV9DjMk17/dHwvpLs4QH8WME5jwYGkdIup5swgCcoziiLcr
PQX1IjX0jZ+a5MImyOTaWzC9Sqstn5gd12k5doFCugIKrLBjR6+kEzhULoCN/2qY9KG4YFxCppg9
ys4lkEVKCsbEjHNffn+bbk/anm6dhhTlZsXoUWjIv0XnU/YczXLz6PkkRbMvJ6Xj9qHggSONaxgH
JN3dLzgnWHW5IP1O9iMFE2CTSEVed9ijVKbSCCOZiYwQ+CxEjhyid2ZYWtZemmPgQ6cqrlcQEtKN
ZQZipl7Xc9FhlwiLH4Y7jIPO6hYPEV7kfrDm2RaoPUGpbOhDVTcPA5Xr+Ebo1wGI5S0HGTQo7PWT
g78YK9wE/tbT3hA51wIj+3Ow4fENcbcTCj7zjmWXo2t6nIWK+w3/77YPl2XzFzjWNuC+u+0vHtXc
UAcA8wvDRgs6bU90OHHZt5zOYI91M+E2zNs1u/KZx/MWjzr3Bj52ig8PsaUXL1DJarOaRc3erP+3
S7wrLEWDM4j5OHrhR2S7a3PHBKY6rmXOA+cyyCsOlhxMKFI/W9pe89evNmjCL4Pr/tGygsWfyJfy
k3WMebLn9Bdgqn6O+hb0svbMSQN5rDdokC3rdkNaeA8SymfSKufIKlnyYeqj2IAf6X8/+pzxNz+2
AqGSz7tRfxTfJplzfPuZnHcfWwuJCvns7SqH507SPodNXY8KLrAiPxAthRf8iAbiM1ekzs2YMMjY
XnyeuA12BO2X6s9XTVxtmxnvlLKRdsfxhTaR6BpSZ++7Dt1N7REg24Se8N05RVxK+6il+DM7yeYY
vL28kVeZuk77VJxGyeolNhHoErZJo+C2y8FH3bzDn/kCtS1ehAZKKI60KQsmpqgUfOMrKtVH0CIz
hY7Xozhc6Ncto/r8p9vzeYB50CDw53I2CQROgom5Xm/8w+5Pr6c6u+3saw43UgThAlrJcen7mvdX
5FQ8NQWsFmWHwFVC1sADNM8AFX8usC0jlf8K+6O4FMilnuP3mbuI/P7fo9l8u8r6ibmHkX9LKH0p
rX05ShwN/Wrna1WQJo1pznn39dTSARMk43FymN1GJ6rhIOUFTZGhtDAXME9qebFirHiQL7hg9uzH
K34kIzVlSAxhMb2WF0TiYVhwyaO6b2t1l3MZLJls4jGUkNXdLRusdRbzy9eVo0YooBSsu5oxTxK7
dn8zC5PneHLffPbaFHxWznDtKUpBKWjlHCFOJs0x8EYK4I/N36L9PNqU8g2CUzN111mvs/BQ965R
WJS3HIsmDabTl9UY6w54KLcUtgf6nxqmCrQojrd3oV4i0YpBpaS6BYHzyRhXpcEVFkfAHgOMl6pv
el4tfyLoUr3cMfLpQBNJBim8WgZHsijhG49gYzCtIu/wMveILerpcXkTCKHK2dDNqUbQWalUuq/a
JXr9xiwRrn3W8IxcT/zkQWyvMXUbJNCF2BgUuQbAz4W02PZGmT9EE/lJB4JBQen4hlMjPKMXEdQB
yxAD5TwCIMnBskBrdjhRMBntwR4dSQEk3n6618i9GUJSOTtGKinM1u047QUF48YbeJMUxvGQQ59T
H1+FdqcyWstao15stC9H1oa74VjhNmnGk8rhJyTby14p2X0Ip1+XoqTL7i+jLjC8J4lnkRC16oGX
33MlKuPJuUGrpYDiY5XdnA9m2fGdn3qu8eltDoIFFqk4kHpR5McXv4YfdvC1KxQaGNknwlc725Nl
jd4n+L9VEofzXhWX/jk9IWZeM/3A9i3bPk9Ix2zBMWL53U+qjjweZXMrQxggirSf7v5cPFV4dBxN
s0nNIM78d9KJ3cbR8fEpcCoQD9QdR3/FO4bnwua84wlEMA1iW+IH+/X8y3NaSMQ47HqOwi2rokEo
Nf/cnFyKXhgBNXyq5lK7/Lavkpyyz//3IwT8k8Hk3JrF7U5Vq//cKyK1ixrf1fMtjbazs9m4tLJt
ADO8yl7xExzEqm1Jxtn1jphvXGw54mPwNeMPcqgvZr8caJR7b5zifJg52rv5Lg83n0RHBAEL6RVY
AOMS23f+IkIboDzBBJgIjXB5sgVXyV+qDKl7UswEjmtHJo8ZE/IKzTMz9cEPgCzutC1e86zY5qSW
L21ebcoWN9ew9239hbMPAsELjqKc5jUFcN18GEv6Jj0HmYX1Rg8P7B5Ys2C7mbgCDwQdwL/JCKxg
pEsz+fcYe8fNIwo4Mql1/aSxukxXPqbD52LlpckubiprmdkdqlvEmDBTl66GERRDos8XhnwXyiyA
ZPNo1hbctSblUoDrodx8nJ9+I63Uafg/pK2TLChd+y2rMZxLkzF0NtDGgu5ScxWJ/I06Ui5NfpLT
JNm3GRtixTeglzYLe3nzoZpQxCKS5/SjCDZp8B/sF+Sqa8VSeb0D9PA3wReYjRddwGhyO3z9sXU9
DxGIn2KATDVIjXcyrW3QxCiXF7aM8CnwNztr2+78QuDAg8iwDYOWfNmlbUNgq8md2gvK49QDoiAf
0y7zJiA8EEsHkpaxNfRDaQNkmWAIxRC/Lq5N4u7xA3CMsKJ8YSTY+3p3NMMwvpfVgucY/PqaojLx
XiiMHo3noxS1VGt/GxEZ+bA/wtLoHOy0Wr7MCM21E3+yec9pKxPz8z55SMqllFAZoMS8kua3tIcw
0dvm4V4TC4JtngFdY6UTHUGbgLNlYTsahHhfvesJ00Ms6TxIUh3kN3gVPi6srPwJz5B7iD7bi1XQ
cLyHDvE5AHEpcLRROFaOd/o1wvI/cA8/3x/Lw54bmqOCyyjbO6nWImUIYCTMN1nxYuWPpZdsjR0i
O0vNf4CwKFbRL9BlCtVUSZFDjtz2ClCsRtEaaEA4YbnU+yV7ueaTcXr/Xazgb+IbETROnr45KFRn
n3bcKxB0Z6Vsk0vTE8CdVvLoSKodfvYUCgjfApvPfAskiJqHDYTdEVtvFVVudLwb/B/TEJgXgf0R
BgG/SPmuT42pkwfNQ/794ItJ6P3IaovrA6PdiXkjOrI3alHsaKPrp5SDf8NWqos7OU3vtVwOhnCW
xIwP4TiNOryINzXFP8i1Bv0qXdl2M1xySVXGYcN4KYY4Rv4RIS7XZn+X1/8bl/cHuxo//C+8CwdC
Mst7jYtX/qUE2hLHbjCxac1w3T/VIgy5yTGIoL00JO8pbAo+VuUdbXFfT+SvY3qyLuYNRJv3FROK
fxyqLYI5y0ufbDHsMvcaEvdHxF4/GnU2d/OoNCqDatfaP2jWX3U4YAbd/aLwLg95K/02Vkpc4gz5
ncOPwieHQtTdO6WPTVncK5ORFUp218iLUlPomCJo173mNDxbqa+iXLZ89Dx0Wbze8/WTXl89lmf0
TJyu59Fk8mzykLoKuWAJr7PurWpC2fD9JGAHtsSC0l6RB5dMmnRnf1zsD2p/pknmeWdWofUh2Yw7
P2UDDV8GSkxBASbEeoB5pHGcBgiDwr5dazC55V4J42s4iNB0X10sEQtJ0oBrh8MQ2NyItDjpU0C0
nhKg89t19AbbqJOoljY4B/ktSHRFHbsorRfBOmbFKQdEJx5g4OYuT4IDVTaL0YtwU1TTb+eoUdTl
KYkLqYTBAb/kqHmm0GEMlGDUzkhtiId+0eVMDWWALLnij6sT8P8LhngxH7Xv/rcUqzdW5yg2zaG6
4z7E117GqmBxUjJ8rC+K2zCWDPXhzMIVqBWsk/3GtpYM4JH9Kblluko5bJbnRb2gTabV6oAylrRy
NCOH/5ZtPZbgQGp0QJmuR8LKFpkPASuxHaB3QNRzwyGHUN1hIvruYoWPc+tmcHnjjjfMU9fpajsl
/8XtUwGmlUjSiiGj73Y+iLnATJZuQHMZ4IuCXcQQ63an2c6Qr8Hmc6c+QWgmpyQyURISYd+1v6v4
vT8DC5BQC9mKhi26R8b5z7FjsS+5jViiDEXQYezPkivxEbkjjq5alp2WDCtN5GZj5KJlmQumsS8t
MVOPqg2Kn55yTP69TpxNwueIB/gFXMr0ISAqGgcKY7i54rGCP4KLDBlCdTU6Gbx0kIa9GoBp5I4R
qS1D7WMUIDvtTuTcJ+lZUmfloV3SBfhScdUYgCvHFdH4dM4+P6svLX5QWQnGTXixXqZvSfx6B9oY
BrjU+OeeurwZm5ujby4dmGMXlle2FKyYOZQEahuQHv3nt/lh4kw8ieIEaANNTxYzlEvYxjPgmdUe
YdrK3SL3jpPR8aTjerqkyvIptVofoJ7RaapKZYmKT7e6FlwC2FZcujfd43RAk3oY1glhd0KD5uYH
/8NKn1Qa3HziIC4ZAMKWL2+01Yh5wlZlbnQ/W7nXsHovZM45grXOFxyYX1sY0Q2ZgZfxh503rsL9
5aHr7906M6aiYKzZCvHq/RE7tzl4F2ZA3tyh0bLWIKHywATs4RsBo0aq6NF4KkHxofAH+23pqK4b
cj39gtj9ghnuip2YpXGFLrdwe32YEHEN/OQRa/zCqNUzhtGYkiBniXS3mzDqGHdf4gVkf7rEXs5k
JWgti7wIWbqGWkWSQSWvWuHTeBbgeW9EktVBJUXl/JuCbZaJEBcPWOQYkhIR3TK0twKuisrYlpyd
F6gTQyzhqtBjDo+/pwhe986QIyxU5PIXu+a/Q8Kzu03ZsZF4SXvI5H2FJAJzdu9oceTcPHjjdq8f
+YfgxFkNFfFChVAAgNJISZcboFeLhhXTW5+wIaEu9thSBtwZKO5E4qNotSXDuQ93VpRnUZhcrvFG
Ctq2bUpPta4+IMILhHJ6EC+BPcoIIwOBtdPwf4ePww2p01cas08hirAnegxZmFdhKqNVPsDZ0RAI
BB+KOeOydDg9IDijcZ7VI2V8129DvQ0cCpy7Zjsv1mPSIVwaip26Opcbvft2ejqzzS+gCKeN3WC9
Gj4m5LWTXF2y9xtIo4x/QKxf5lOeKFUhpz51OBVnH9hzjt0zSejq0aHT8tMGF1Q9In0Qs+khP1RL
o4Qo0BwRvkBPgtkJg0ebYIzFje8XS215rUa79HSfutxTv/0WJXx2EJ3lcHBqK3lJiiKuE9KPGVTT
2dmcYy8T8LG+VWJl+gyrzO1HMZEV7+qFvMUlaOmnq/HesSHQrvuOa9QV5WGpXi3ViWfTflFhjJbL
WlE2TLfAcDdDR7Pk2FCehlFxFBIS17KKXWrWeY0WX4OFZoz76SxJmQ+mtInH55sicwfMQFiNK0KD
BhCakr45SqnoosU4opy+k7l7F06Whx3lQDNBDLaIz5ujZgN6s/Ia87XiGrs7q5KSECK4uRgaJ61G
hAv+gE3i1ppB3rvCwktSyqAQn7Pb5YQHlYq4RB3iBtYIS6pk6DBqmy56UvY0bFCvEbeg6RM5M6pq
c/pQpxLjbAEOUZSK6DRFo2g7f9Y8GAsFgKjae6NoJ5thJCrGyN60zJC+ntGWEOnFvQB27ahY5vsX
YlZXbCUzgq7vie3OuSQwwqbjrwHqTPxiJ7a792LdmePXYUOYSk0FZzhyIUiDmoQITtrgDxhghT8u
GHoerOZLfbmsAcTju7lcts4As4CTNSQ3utPdis5W4GPoncK43k7OZbXEgTmkiNc0+o31tw3UbxUP
5FodjZy4wXRtdQ5mvenXZzHHe1tcX59Ok0/32ECaCSmEDiabevQn+XtfNhFXcOWUvSN7RO6leWhm
Muqcht6gzBIsGcVykDJxcaTJ1MoMh/9r7ynz0+TKDyx5DZKttQ+cu8CTyxmvxscF2XVpfNiHM994
3KtD/7VZhiilqli77j5oyMGM3Dncc+SYG8xsAQMlDULeoyFsy//0ldk/942HwUvD4GezovJRxKSv
pa9eBiB8XItMG+7pg/huxxbLAyYxRwwmzDsKout8WoGPwL9Jyp7VmeirzuutbcGk5QtDAKTXxano
wYrSaF1Y4Yl0w2LDmYkZHPQUZutsnY2FcxqoJ85rVOMnGK5a/EM29vmtAaYHrDWczR9AUZVz5g6r
opw6vfJRIl4oiyXua1YjXikLuz0DHVJHBZKOtkIVq6hfeUqXu2tuQlAnFXtI20eUKxcTdpoGBwmn
F5ZHpDMLiFojM24RTpxfu4kDt1qSxCk5H/mpt54IbOT0i2XXdnQSoHe0Xxz6GFlU15RqYROs9C2E
Xgcoh9zKg1AS1pXts/RHUb17XGwVRJINPu9Rfw34WJv4SqVJG0NlhcNhNrLonyII1+V55EYsEAoy
XABIOvWF9Bk/sneMkXiSQYiIcS6kxuQkoW86e4qDKJUgGfywCrKoOmHFSlX+8Y/Tl19omrqHqlyf
EGcqYSkz3O9JLygVgSkNZlxKRZ2p93DarzHyU6K5JDKDVLtyeNMBMnZa5oJrIaupI1TY9F2qyeV1
92awTy2NSxBULS6iXm3Knm3jZHLwC26e2SraN11ANJkzWIui39+MPi9+onFHQH0Yk2KMq0Jvk+Oq
ClMFJlw1khE8qBmWiI8v/aXjJiC9O6ddzSS+jiIvcsKppDIBqQbwyg2y6O6qMPrtY4ivp/PHBFLQ
c4PNOYsfHx9UNGKbYJLZi8K70zxAhVBKHfUoCVH1Fuko2x88pp2r1W6Lfp5FfOj77MuMwMewBwSG
n+aLuECA4ZHLFybRQk/UV/mjD3nS+xsJ6BzjV4o1zPmR7VHImzRelyEnQYjOn/pU7yXs0vR5OIKQ
+gEvnth9RQfXvV2xy8kg6WdifwGkUpw14KjPpOl0KnYXkY7uUcrTHbgSorAD+Caiz5T0PDpSwbaf
CqCc54wcyTiewLyFdfHnRkdD3UvrM8Wm55KiG5hfs31e8rIrK1PEIqw7Sgo8ouvh/VWSyP4w11R0
zcDqxGoqSNm+1ODm3KYbGDTpkoift2HRezLETUfBkCH44FUxFkPB55MyD434XnaXQfD709TjDlu/
5XOiDsr4FBnLlPASOSrksRADqTVMQMXJvcA1KFd2LFgrqxbS1eBJOj0lU1fCvNP0SJ595muELRbc
r3WL31pLeH2TqhM2Q0AcShmayf7cqM4QDe8WgJvW1ZACc2C2T4C843LbqsO7P/sBTooxt8D1WY9p
zu1TrINUmWoKly4dk5hwjQg+OnM3Iy461el1yJ+va+S60tG/R7eV3Suf3rnSJUNv+mYhof2SQqRz
FHFD3wloWGKvd3LATSJKxx+KQ3O8cHXU+J0y4zv3h1TRDexhY9/T6cOLGxuBnyY9v0a3dLBTJQxb
UOWKJJFcvYA+udZmt9qjqufzC90q44vkxA3HrhAZT6YF9DNf6mX7DnrNgu41kCyQ2CCJMsfbbWX5
J9oamGyFVb3AxFv2clXzX8Gp+zQgcAQomkrXjJrlVKepR4TqajBL8BfgL5kZEiuzMNCV2Xef8yGr
/BhpdkPDZNwYYQQbnhJmyfau0APkkVaA+8v3CuDqn7XP9EwXYzwNoMCNN45mbaBrsd6q500uI7qD
UvnCPy+lj5tAJM4++gZXKov1NA2lVuS0Eo8LkuaMmzgaPj4XP1Oalq+prsfGr2LUs/qWFiZnidHq
LD2zkHjFFanoaKc2DwhrUYcLKQzK+3En8wF/2MLsRPe4H3MMKoOE0qzyxFFvB+LYbEthvpPUtNSB
YkoI17aknhSAryWBgXvi3O3kiqXGhwXxuNmCrgnGWFVDSsUZ02IQssMh6SGmRTaPgMeVqCyha/PQ
puIha4LaiGeXP/tcxiR5+UvotZZBV9lyHsKMGqaqqZiYeZ2hI69gWnIoGAjGg2aA0r0uEvLC/Lrh
/QKD6YqhcP4I2P49LoKryIotPCMbApJJ1WFuIXInEnKnj9ydajq55wGtjyNyLm8m5MO8VpWQDiYd
HnuHqbKQ/cSMtvwiFHdOMk0bmZuZ6bKpDYmEgZSIID5LKAK+SAxhpNEvWkiVtl2v41IVjeD5S75B
FuwrsQkfh9rinx/lBB9uYFKD7lsC2aPn3vmmBSpJzjEp+6o7LqaPEtxYhEYRwAxHuSY1jUCjT4t8
p10M6ULX8azMbxMwuDg/4NQ62PBTcmBI10Jx4ubaymfKNOMp+PgfmYgJfaxCALbXrCFsrRbv38uA
xiOjqc1/dNrXiKuniul7RDyiUhrTrWVAyG1lC6O3NvxDLCMVowxCcFgKBqISmwhLrcQJU9r2A/oI
NSvhomRo6kPGG8n7X6KehXF2HRzgncbBjE04BhBsWEZWJP9JwBay939TnpsuBceEMvdto74vbWuX
lWImH0a4+14FZDlVwW7XiloLEPgyahMueO3Qohb1x6i6tj1wodB8e0u5rIn2IniyC/LVIW9+BSXU
D/RIN3rSyOMT8yawy+Hwh/eleeuxOflIJuAOrZ+PTC2RdC/5vFj5YDCfw38yh8iu4dueFhvV5pU5
Rdbz8W8iZkgLYEXq6R9WiLnHdN6fGuBTldbG5D72Hpq59aimBT93KGCmONQ6tNIE1//oWY5FTXpR
VpEEoV313uPK2Ulqn6r45LkeMVofIgz01rcWfmw8m8ZnWni6ybOYFKWYlvHI0FaXqfF8NhROPtoZ
MznWRYdaeJdT7+o5u2JUGkkn7oZ1WQroBjKmXNqi19M7wpI6+2Kjz/G3pM2np8vSVPJNDnJQMtTP
/NEFLif7NTeoQFVKOEZsA/ac9omGpof0AB3d8G06lgujOzxk2MF3iT3XPJAn4RvemHq6D6Z4qUct
SqXk7ztVF1AxJTFd+BBN4RE9SFpsJxpc8JvPGKRmHFPYcSZ6CzJYFwDtz+ceGF/9A/Mp17Ra1OJ+
UpvfRmVSSDdLEGJr3kVvzB9qfKezxuX3cVydx+u3x7luEC+fGgI9s2mlihUun2AktLex1fJSPgZG
uzqznAHgbfrHgVCtdIR1gQJNwsW4zJcgtFlMmct7ozy6I1wJnQ0sO315g5CyXyBUPdEkIzO/c5tl
A6hjcfjWDgh8Xxkusn8amriL3RW7gAgf2EmrpL0rZPV16Cao4rc7zrF2+nW1gtcDw5eXZ298GH0j
uJejYanf5u20ij9FaUsIrZVaiki1yMrXBZ5n8RgjsJU3uahGoR2tS7VzI0A6UcV+OF85DMUfl7dX
JQ+/Zd+hAjhg6esHG6E+vgtX3IFiLmVeW7OxzPBB6NX2VJmnEUwFsmNTJDeJXqj1ZU2oqmdakay/
3MVt8pPD5n5LeM/KdmxVIDgoM0bYmozfb3V1G6LqU1IdBFEbEl7q4nJ6GSXO2gnQooZxZQ4IVSdD
ijgq8bJOfFtt5e14ot5yZGzgLklDH0aiEV8BgWrpQe35c/mCggRiP1txJR6Lg/2Ou0hkM7KLvMML
jYb1RYtY1QgYRrtp+NWDHgWNUjGLvIZJ/ZnwFQd70kD82TLWlTEZOVKef7Ooq5/0YzdiH4mJqWdh
D7pdhZg686H0XyeztR+7SSowEgPfnCJtRZ+QD0GEjseZyWfNNkTc2UiF27Cyl4RduCjVzv6O78Rd
QIevd6quOZ4fM7Bfq9RNe6ZwA5MyvTcPEbaUGgDA2qZX9c5EvS1ok2vg6/a3n5s6G993nozBKtJH
d0M2PTlwECPq7ezMXWd/qy0+a+P/T89YEUt4TPnZg/MhSzinMQPnPCfuQv0iJ7GH+S3s+YMCrnPF
XLVMpAEYOGSFIkhaCrCJSRX250hg5Kwze5oTf15Gw6JiSIIjnyeKAX9U0SdHvljLkLxFLVfvN5K1
yJh+rniL3dhdm5dAcwaywKOKL+AnEbyJQXJxD3D6tIbMomLUtragMpIBZdOFIJKABSHb7Io/rNjd
kKGD5Txj41Tbs3J/ovsdtwbn2gDCbfNHNT/pv+624vo50wWjnZNzuObkMOhGoFRKeGMKbmiHzZHX
ePzWMTqwwLOhyMSsW0RWmYcVvakpbNWOtKokBw15uP0MvgTiV8kHnnuUrKt1OknJ4OXS22FjsAD6
nJH8p+h+zyeyX35qA6kjux/Ncs/yoOByU1kXnRbm2V8vK0JVDTH2wRfHMTcKUgTL2AZDqEsnJdS4
vzGpFXJny7HIXY+PewuTiwMKrxECXP5Xr+5TbTf6xycAc1Fi0hpTgEGsvcfFzjytTCn5raiKNiL3
Ahwb2WGYrZ4jeTchh64QuC5aYVSxJLYMS7hNo6Sw4W9H/203O4vQgq8GuQuHDkHuQgImA7P0AiEU
7rSlBTWrylYgh1TS70rpmr7/tNCFnyQuNZ/eyuguCUGpn6v16ODzCwvw03w67EZIq+s/PImrRQG0
fnv4b4SMuxNq68wLp6j3qxTLIQiQ2Gop7BPFIOTCGb3fw+N1W6NviyWYFVxKC6QE2q3e68XofQ7v
Kr6MNAF46CH5zdpig6CpOMxAE89Jed5XjUO9bZZ066topR0W6/LCuM7dlQHId3uNjscvReQmmQec
foGjh8KJqjOxHDRPlFBeABsARSKarkCu29C/nIt5vBKQGEYUQjz77Dgb0UfuoOUoN+aYMNQDz0B9
0X8L+tYsu1eapd0YNqQox+ZVZ46TbpVShXU9NE92StlqSIyANR4quNO/SgHRZ3nF6QyzkVvA4NoO
rzcorfKQfq+G8nnzi7NEpPeUpZ5W4pAlYinSdCtA+K9UZY4tObCh+BplCJ8908xQo1gRGR/xhyar
Kn6eAHWa2G/cCtEc0Zrt3wmED6P2i4CXxXvr8iPipFV9RftfcgrhHL/P0Vz+HT3ZDiSRaSxnEPKg
EpuQ9tZ6o0Iv168sGQqpohMMizVcdhD+AAhBLLw0TcFl8leRdQ2OmrEZ1/1LSzZvfAmA6NqsEQwK
PFtVmOEsH6uGGrNHGYnkAaT/yCAZ/vpwONJ0zD4HqjZgFGF+Uv+3BFtxefPO2TB5k0NFlGAC4lcv
Pf6aJHhJdL4745pct8sQ9XnQ373d9dFzKM1Hm6pGEyqlCPW0G0poIB8fsX8KlweAPBMQjVGcWRyF
N96mdCXEZ7OzaimnnwFW2upUBEhHsLRwD8RRFN5YwCCWhqqYD002b3Dwa3Ob2RoW4baxBmVv+rLj
gjTf4GFNrEzbOraIrnlxWTCEmkfmjmEVS0o/xMLujILX9u3mnmCXfeHbaitec6mPj10yp4VGJIhS
eoGuKLFcTwSEPfSqr0QLoG1q9Di/Vobx/msIVuw7YPMKMXyIHsEbkKEszLkwMf06TFHMMPEHz3pC
IjVvShJEwEUonyC4hNVkxR5wmYemo6spUNfx9IpnYRib+BnUgZYVq7hFF8kPNiuYmBnjFe+VSYoz
824hty5lEu8nhjgXIrAkUZMBTus6JusSSNJYj9Pp9pqPl2/LXtTlSFbtjlDSXegriBLWe7ND8WYV
r4tbf4joqDyZKylkKSFgSf8413PdSwagneuXWstzzW+BqTLXWVpfpZSsA0St3WIa1Y/BcNZopLaU
qq9JxAwYPkuXuTCLHndIosvQbuIpjiYKeRqdWcgB5SUq487mD0yDt7Bf4a1GYjehXGzJl1y5FD/1
BSX9O3pRAuxxSAGPkbRGGxemVJM2HNLT8Fc4KAQAfVNSIpO+vdPTn95ND9161vARRhgGy458iH58
7ZkqzSKgp7zjbbJYDf4R4pr+WIBbeqwPJWRaX3feNTG9VQhMl0PBlHorpiP36os/FyEVVob71Iws
hBlShLylxUpgrH+hKyfoEZNkoJZPrKIAQj0EqANVEykzVv+sj3dorgo6ZxeObQ8ViB4NidhGw2Yk
x7r+h25b87z4P2VG2o9dgW6qf73jcaKTqIpGHRDRa1bTWV9i8pOmIn7qJkBWvTSdCBsOTQwvBoLE
IdvNZLdaHoFx1bvWspjStkNNYeb6KtnKjDNO+cxb8BHIipfZFXnFnslpTPGi/xeXXUC2a9hlS3TI
A8Px1qDBEe2/58Xui0zBO5w8LLHW5W+fHLtPBvQzZ5VZpWKUO85owmeUl4cO1fdeyL4D9BHAi24v
AbEYapagwXbypoF7sHXM444dUBfSWPN9KrB/gHkOlQ1/Wvw1Z7dwdXMG9+ZmFKvqPJhjZsRQ1lA3
PK3fyfypqv7j0x2SKhen8GYLdpuHMqMRzR1KxMClRB0GACS+hcPFJhqPHnQbwplbvfXy3S+/QvW2
uXVqQrhqSIKbthypF2AIUyZZps3RzE6kxg8VAuqKZpjyxv9t2EPK3rz1213g8S2oO0eHKr1xWvoV
nE4kzLdZX8dTc1sDvT0SYi2KN1Ngh6WA8ZTSptGs3rqfEiN+IMkYovojO1zOy77CFOguWQmGxcxE
9DiHAgHZqh+MPUCgdPYoqn/JtnEAqrg1Lr9TiydHGskKu6Xjc9CkoX8oqdoDEr0A0AUNVeho6177
Mq2MxK2SoFC1arglawl1+tFbK094Ffa1wwk/1NLbfbtEN8z3GQKhUmTg7Us9ymXJ80/gNRIXxgmo
WCkBeu1WDmT5XAttSgNt5NZ8smsB3SFswUel53JJa8sXn96PN7vosZjM/qtS8nxqhMoFqID/Vlqt
X3PaLUouxuPTP2ZR4ltuQYyrAUEp6ZLJNVgrMc6HtX35K0Q7z1smHuqOTyVjPQgdcjO1YxDvLZFT
J/12OdhHdSYW+aCAps/jy5BG8hjz3V5VoT7TG8mUpVqW3Sv4eGa9tmKfCOCjuDTjQcz20ZLHA8j+
iUJeNzW872/R2wQJ1OoX7ntFH0NICGv35p+Ar7h+3uYSRrV7KC3oiu9U9zzXAlqAuW9NSmHOeHHg
/3pQIgcBCif1QPqw0m2VYYPYU1sFNasW8CxBnCFYqz6e766wvqpaVjaLIn8fLOPIp8Kz2yuBOFgV
21KY7OWu48PC8ocu2mlDPh83QWuPo+rR1k6xqkeW9i8Pd+w2pmc1fIFM/wjKgkzR73Fhv1MT5hpL
Cv1LH8J1715vqvqGHgynx6M08Db2x9S5JLOYFAyghYk7GC8LvrF/jWxZigMDTq/N1dS50hYHWwIS
iQhnkvQmSKaobueLo4ZntQeoAQsH6SM/csNkd23WGwuB82UrEXv3713R/+drBx88LNqmNcvkndvh
tqGxEWAuj2vXvVm2LgtuL0uUXXKSusmHyVQOHTkRSajEVGyaCPFNmqKCz5FtAJAbn8T06IQrITfl
W/Y1dWKBUaAQqaxytwROHd+vBjT7tOpvZhGpXCIJyHmOQTHOdRgJQ9nmPwGdDfaIB9XJzbg4psrq
AtVLctD2THSTK0wsTkusSf96TMxQ3fvyfmX8VNOod4ckFgQHWRkfduZ83JEQXBeH3bQcsHJbfU99
XhMSWeNHhP9Ggcri2FotgcGMuwoRQzcMrRq+x1+p63vDLMsBmwmzuoGvM1fG8Fnw7Pcra23s0YeI
PWeToraEyacIftLSCU1sLAs2Hz5UHuoTNKCuwp2qdF3Qu5ajxtaYZRXKRmDmFBnvbErQQUit9vsg
v22fNf4drBl92XtXOTHny8RCurbI+BFyLueUgDbORhoFc8Rxf7UmyWzaj9o9+jWqpRJKkrnz9ChP
NJHchyX5QKf7Wgg+Su1dh8+XCenMaAAg4wykVuX6m4huJB7ARx+/gt9XKMgnURnAv4r8IuQ7miwW
QEN9vZW//l8gMx/GCFPTxSki2OkVdpS2qIqZ8A6+l6qBuJg/Lth8LvByZIVLuqAD9AzbdwkdMcHe
R8hLQOBd1n86YlDGev7u/+x83YBGKPl+xxtKpCUaLurt2NGYk+JA6f9QtrLXhGr3SeCmcgQ43gkg
Z1KrIhEJjLq0WLzcctjxx+KMlErO92Z1qKhSVa3QMU6BCdOTWEhRcLekaWPiAvho5D2AL5CKZe83
qGGBAAmnnSNYvbO2tnDeidAvWjdrTFkNBL8mzyjpDkpDEa/iCI6WQ62LT285BwmOjCEhN+moksTi
7E0PvKee+XRsuw38/BHRENx8aVGplfGkBO3EvNth5s4hFwhFCMeiwNBrFtGlmQpj/4+68UE2QQLB
nOzVDUEp/tA3PoolDf0Kp0KcJleeNU1KL5SLC5Vt+dnpP58+IYVFEkYiDsaMI5zthNdSWRPm671c
hcfkNFDTdSEM3QscWuGX+94znsGJ4nzMHCn56xnn5em8WdV35xyoZbiYjO6LiMlTLsWcOTLhe686
UPqAuNa8sUwehX4TJRMDANbKhcPUVHtfXRUOl0IwYJv8Hfs0n8LT95+cr7oWeUegsGBR1qMlSnrQ
LrNIesEsPJCyIMxfhpfDDHJSgblv/JMUsWiME4AqIRTMgFhUbaOz42zcUzkS+TyAy45WgJkHdp/p
hT6SpYFYAXOAMgapvXuuX74UcHMqoCwUJfsD6Eg2fLdXyKf3AGXXp/rqkhon0splo5+ZRRKTq4po
qKqW+b5dCKNg+RCuvfFUOcBmSqbbyUMkrDVOnGnl1DCXCG1bRpIIY07UlAhu8QBNaqBjuKi3GHyR
GhMWEOHAyZSR4stReq2aF0r22c4I+8T/22b6xvQUu1SXWDq9bwV0zZY6IDtmvyJyRx2rrHBXcHlD
+cKx/7f5xUnU359P3XfveuxDuMMgq23iLiQs01fu4clcDxxxvSqceUUDXXqjCYvAwrdnD7KA4b5a
PdKf5nuWemM2cQ4On95kF5tqKwvXvCcpwzqe141WsU1WmNfHdb+Uu5oUv0CtLqLGHyfCoVCZ6Exp
YDgJ/EJ3dLpXLhVp3VQXo58gZK2c5ISh8EQermqghRuH4DV/hXnDfP5X1dBWksTOEKnDOrDzdcFK
X7s5DFS0ByXbcbbJBzD9N1WoAWty0ZzKJ8tClQfg3pQtB2zdEZZicxdXb7/4DUs5W7m1wgXNhJNq
TU7sJy3dc4NLgDpiwJBtr/KmdePmjshXD2rOBzDuRBFJGG+qVKPLDjj6Yqg45qUTV345qwZ3KFI9
UWOi7BIo9ZIQPRtc4UrU8jJ4l6ghd+GF1oT+19wWW0p3KnhWkq+09qEWCBvibogQQqmx/X+F1bI/
dGaEgh/RcUYptpetrsjNoxVerOUqOHkWPFQt8Lq6+S4rlZfUkFVbmuM/2AQF8taiWeExfezptuzt
Ghps0K7R50AWgWZ2cfrlaQ93xMJKRiO04Df/Bc0iiy6tEid29jjqtWDu8La/csuE+3b8B06YaHd1
UPVCPH3egN9z2AZutFFBqGB8JHQw1bm84yVglMETNja1VlwINKpA/tXoJC6bji0N/AyxlTHzy0oQ
5uloz2ik0IiGn75T5goXVgSxX1mj/wxOcrVcWiJwI4aMOvosAO2d2RBI/KoDVh52/p0lcR6Fe5D8
FmSRCZ5jl63PBlT6muMu73ISznF/2DW39R8WYRT1SM6ZxlG7A20t9bFF5XGwaZ18Vvud2bl5cgk3
nSteGtLiBQ1ym19PT2TuTiw6qybc7ouQodCIAh1XlFv2OiDdgXm9IY+2f/ib8V3bhOvXU7rnlT3u
RB28jZmDYwLgQVDnZkM9W5LsZdy9VRBYkVfD8be0MdDz/N/whURBJmLQcCHkKN64e/NWwceZ10Aa
wI31R0ENCfBR5kiL0bIe6oBHdoh/cMxe+UwtMeqpLT6ZWSICRmT7NKZhYwseQcA+Ei/q0675JdVU
SkWDXve7Q6uznw5FcGQkSy60pdpy5Hle1jb6KNVfcsh7nCP34VkR6cYFPMuD2+Hx4MxDdR3Wu5FG
u3Jrfyt0YIiP0srsChu2ASpkH6nETBPCJBGbdf6bdwU/PtAFsgfbfWjVu3ONQ55aUhtqrUjxLHTo
O3lZMh3vbglWOLWgI3ntRgaxYFWoz9g/LOKa2EdiOcukE4RyoKMnL3UAU2PZURRsHuAQpX6RN/I+
Cu1xSv0sMj7/UUU5x1MVKaFg0vE5n4ZaBtV0m6ua4n1YKrwWHKn5N6C5nIJiemryjFu64oIpc9+/
dZ4qXJVqQiwBvnp4bhfQn8DIgehgXbl2Fs7Y/mAS2dsxO4CByUkbFROh49WKZIlAG0lOD9eGj6RQ
UfOWoXKTAmIN9jDb6qqTKw/6AAnmbxWqofEvdCsS1YID6XK6oL/Kp6wTAm7l6S5ck17nm7GFQB7R
9RwtCDYYVOuAHLfeeo4D0mL+utyUjlLN/8fiH8QFgfX7E17juz25CXlQxQyxm28ZrRIir86e/Soe
jga3RZfb5FQSziUCDOpsFazyNzzU9bXOsVfl08tdMJ9BHItWQaZz8YMfhSr8SXszWDPmtrgoo3EE
uTGpYrk0lbUgi73UE+g+WQwDVbq2ZMngrHZBRAKojkjV7aR4zm/MNTLZkBUgE29SpIE5o4psuNou
uRYD12eSqSB3MNXhqU3ec6RKUx9R4YfrMshjPX3C1ZK5jY5/76guOMCLH/h2GenrFDL86DcbZ5pC
O9qTArGpc8WJlYjYJ92HNFh75FxlT0xgEqX45lJ9r1cEUW7bO5CwHs/U+lNZp3ciOHf1rDf5k7KD
mlBhrSrL5cFLFkph18+tFzxGsJcbV95Cy4pouGZlDhtY+i7Asqqgo3WyVNMOSptUCl+m3aOLVSXD
3uzbOQhDI89bMp0xxAY1VtHXcogOMf8yEm5nJPzWVeBHYrV0idS2j5aDuJOl9qOJTkuJ0rRZfaCA
v9BTHnR3o2oWNNRv4PRp9/BMpAShRLCEEDCR8Aui4tz+VGvYtW4v/waFPPPESTv5hnNVWoEy7/CX
+mZ8uKUXSR1K0iy+zlnfpNxSgXk9PAcWgdQn7nlV1MIy7KmJaT4GbAoSy0NU0oWCgGz4AWL2hipg
lY9R0yeI552owpyRVvjJXYL1U0N5UV/7UxI/pIRNfvdzTe6LlrAvVNdK1UCR9k6Xwjs2GNFR/zA5
S0QJcRfrn6zfsTGorCGnWnQWliUgAhWafnt6PNVop8S7tjkTtaXtLdvO9fG6E1+ISwzHF+xZl23+
Cfu1Bj+7IGwuQnaaH2QAwTMZxjQKIPJOEZld15ea1eWIhJlt3M2UeVbI9OfY/Tbn2cKrzz8bQp+c
s3WyV7nAJgf/uu+yJ9oJ+L/zpQ/YDLkRh/iYui+u/6/Rrpmta+niT9/+zUgySaMmaubkDzQ9kdKH
N1X6ZWnTKtZr/udrGvMe0LBVF1HWoJDTCU6k3GQeepvHDomTQNcUUsUIqfxbdKDlTvf1xecCtW5C
k3K75jRn/aL7XKFhO+nC4l27jrDfVl3ifDFylpbjdKniEpag0cJFJ5x6jNf1KVkcMS0Kv+zpj06k
LFg0xUARrMymJ7eUMTyRAxdYWKJy248Z1I5vIzJr3Z60Rv6PV41lGTi4d3CGvnRBqbn/s/Ngjqys
FFHitK4HvO1nUh+w2Knp7FsCNE3+f2j3hGK6WCRI56BOMa/6zqwLZZjbZqP2+XxhbAeSqIrpbSbJ
8eYjqY4L9UdImQAwjglHyOfEfGwsHdroy1ipaRQPnoxYIdzBmk0QS962FXTr24TrFn8K0XCa+Xki
D/UjbMuOGT7CJwMMj/7/z+OGoMc1D9N0bv6biDjalF6MgXeU+BOhLbbRMc+zj/4dT0U7ZHAmen/O
IUpMp4iKc86MvCEKuDk/ohVYwGNAiNE//qAJ/fkSAieldHojAwi5g058rDa6viuZidzObWJmWfDD
b46Nq2GOmbpFZWYp23K0rjytmFcaggKYQH8n1qUDq52tXVq1TSftDRtMJONrHvYOEZUq1XaZdiXn
K0qdhFtaexjAe5V946TL4KClis/e8uGxSU/LHVFPgzsId5m61paDo/drzVOalzl42IS4p+RpMly7
eMRfmzFXV4oUwCR7gJWoyFZmPg9AGbPln7qq4Pxh7hdwyAzp67qsOhUdmCc6dvf7r1WsnwqLtbYL
WCDcEC8z3e/R6vJ9jbxP2AmOHlSdf6RLJEnFtHd8XSEpPFPICiOeGzAJ9jGSbNMru7660GsmGmz1
AW9LRduzQ+Zp41PUe01p1EiMZ3dxt/vqSxjudDbLlqRob5W77EBp4ujIe6qoMYqbQDglSZaEEm7X
bF2zfyg9R/ro+QG+EtwPqw0fFQJ18Cm/uanGAEsM56/jiUvG7/OJesfzTYSxjSUru4mYzQQgV2l+
JvakqOgz26iEdkR91027Km4UPnG11HuDp54A8vnswDn+c6nUZzP9H0n3YHzkAzLSAd+5+kXXt61z
w/Qgu3TZPmfZPXyBv+qVTo6LDPA5YxfoKczOYrqlD59UpBhrcAOgVM9ZEgyTtZcex/5415BRgLRo
0APhrQXsHimIm+SouVUHxYikmDGnQhB/cbyJfXpCkvGwJfxaAlFE38JmcO8MEtSt0xKJUDg8MwtN
EfL4JN3tGXTVk9N7mLBUbhxmOxZ2PpxefpSCBDgFltM8B9xkglsEP4cAxYfDN4WLaSZecCn3PvXb
7Ufg/slpsCBqJkwNBieFoHOK1itVm0NBGV6n5FaatjkU1NZ3Pch4suZ2R3xwb+YHHLKIOzwi6lpC
emE9K+ZAa/1HjJOjy/SvoCaf8Vyg6oLjwn6pI2yNcOu/zDQGCOQSfeoEWpC0LMSuEA5NUmWjHJ3N
tFuUPLVmf6KPrgsmPI0AgKUijcL9IYtohAurHUE0PSWO/OOqtBu36ieovccwq7HzlJLrsVlllH2+
yl23OeGcxQ/hUs8hun3U3lNWp721kz7V0CqPr2NXfq2mDsiahTAWYlej6K0ssTmsqDWnZNocDbRM
Z5Zqr+dlCQsAQynCYh7/j4LFGMaEGttWC96XI/50s4KYGctC386vHI2IXOTWK416W7BVTuBjHtsx
noQsK9OSOpGZRCXnm2liK+dHzeomDbRy5AySz1tojlk2VJsvoFWoff/4U4cZTCt8+5gko3IBsaS8
mZFZjUzPx7JTAwvEolFswPr+FXXvmZdeNbysducJNd+RPyylN1Vh85mK+KvduB+j7M9N+Lnp4BM/
dvAMVrZSbszsfy6npqHHuIArBMWe6vXBik/bL5GrcLLn0mGP7voE97BlRXV+vUwHcsxHYp0izV0m
DDeInR744+7MuefbJO8jIT2Ho0zNgnsZ8xREMKkxZUdGx1lXKmw9+U+V0QYBDv4GLoaMEFl/ZMLC
Wk4SWjnl7FYxHc+En+c6VMQMaX0J+2Q+Bw1uCzyPBs7u2tFtlxlOYCvsiXI/T4R6Sq5ZIPURmT3y
cL3ySfL7MYokWoWOpznQ4jk/HVT5cr69aGJId60mH6VgnLz8VgzBlQnl44cyBD4s97PjbfW2S2Uc
Tz23zT++JBVcuAhSy98V0dNkpyGu1NUXTBX4KLLq3aDIBeC2awZ/cfnd1ZlmWGdKE/JVKoZLvNhz
VrmzcEhvC4rQdqwsMNQPuKEIw1xgWmkxym+kCQMW9ioOqyWhq4TKzNOk0lPCazJHQJSumCmaZFli
GD56SoUzJ3xVg1a6e9B49qk/h6+BLoojPa8XJRYM2euVJ4kNNE3IXa/bzv/EIZ+RS9bblURXADAT
PekHRu43TYtgP6uy0/kkjM0z6u7XG0adTbOrNkEN6BAIMgxqSrqGK7GdrD+8R2kAcm9nDprqY8NM
G5kXBXXUXmDkriiq8Jm/jpkTbV3oZNrMIsF4AKM6JpBBDFP0NfcmqVDRBB45+dhlNHtyabcULWPS
GX6wyRW6x/0zHNzTZtIwOsei2cBnjHay0hwyyU1OnYxS8T0j6T9R58iDZXqaiVgqJsv7rSo2Tr8t
5pNRxZKSjbovCB9zSTIL2hBhUPqOncDXiXeZi76JHpBCv8+1TqZNpFT2vVw+2ZeQAGR7cV+DZUD2
rmstrGgi2QPiORygcZNG/caScI+Mp1MtDsPv4snWOmlXLGZ3lCBh/Y0ZJcQTPQ5sanCUfUjqvFv4
TEetsdWXGgdsHUVE148iD6ttzUqzTnVfGQpxJYasFXWzbRl4fDKbeIcpmV4PxW7qS1YhnttGW/15
RSeWhBPoVfcHXOu1uaUb8Lo+hQxYiLzAJQlg3h9ZGN7z35yDGZXG462aUjs8HJlUZqpQfhvd1SPs
NADMs9+OP8H5B9DqeqApxYTtIHXS5FEeUd0aIoF2iZHVw0x05Oi/Iw3KRrN7UEq8h3rEKhcaUKs2
qFNYwouHpt/D5IIeVfXJIDJJY2XnhoY280ick1U7gk9UBpxXzHpkAthy4hRpDa5GC1CRY+k0Mrfe
FCil6dEi38vSn2YPBdWAU/6pqZrBKv0toL5eahybGoYB4+I/6SWoFwwHMyO5/A0MwQdnOIBlrOGL
/OAK9IlvNRzAi+mXPwwv148uOQUlM3ol/i4msZnPMRYLUYnILO7WitaRpcQrVUhemrETFtZ6Q8sr
SsGBvf3LYNxU5uejt9uqr2Zl0OJe89xrkpTr/u0drCckV187tjf51u1TXE6RwpMZrZNxtOTzGHE5
ZnMImIes/mabuYBWd6aA//o++9bqDvk+yswKSgVtTsHPyTIAsUffwOdzKsrf+W7fDQHOM7J0Q35n
jN5EcPeES66Ci4f2qbdKUgEkOcRVSB1CQniSulWEx6zlBS5KzwlCXpCVOAs0382dZXWpYALAogUU
dqbs0OSC3THcx/K4HI9+Xq4pxBnK0x/vUrfqOEj8mDnmk+nvJx5BG6NMl9Zfr+lKtSbQcyB5rklS
xJFrlFtKPUmz6+EIYll6fpXjgFfNWoneqnWCVB4XRcEVY7SH9fWkz1SmKmodE22UBrqmuMrX7n7W
+oFLoY0K6cT1WfcR367CDUIq70U36AJjrSuILZSQHXZQqtEVLFnRChRWQ80vqKGx6xQlRORTAmQ3
TcbcFBAm2uPdo1VhTjt9EzDPcXDAeLsQSoE2pL0jf7Mwd+ikiyHW9zZ21UPoAY04NsMFb/0OsTjx
FEA7caLFj4BhagrvrlOKWfAENP3wRPuRJV4pwjyjWL+baZfxFqmISV8R8mEx6CX6e9PkvdcH9MqK
Q8TYaYaSrfzbQqq9vExbDi3ElzRVGo04IEg/OrJ19JrpNyusatmvkvOzk3TiMeYWe/2zpiRz80mh
+FXGHb9NfDB7VJv3YcK4oYC7xOvD10UDIZZHa++j97RBGquiM9d2mWnnbxEYxIruh12kAcXa5EoI
cT5Bfz6E5vlBH1leexoUAu/R2lwqsrWPc+WEldG3vWQA+IGX9vPPyQwyH4cjUK+RCRF+JIk5fQo2
MVeyLcLgtp+HsV8/G59fpJWhPDAuM2Z2UluZN5TfupHGBMUfF4exubZLWXLuHT3voob9UiHgypE2
jVRZnQmyChrtJgnfsnpi2ZBBmTVfMpz7J9EsUox+tP2g70EBrPxpIuW7vGpYerJTZdqykiyUq25g
Zn8fOuVlbfA138PPi8PFSgeJpuDKWVC4JuIopMNyQB/fisTMdI7ODy5sAKSLz/L/+c343dq44olE
yxT/GII4BWzvQNsgvIAmcjiC/n1GsoY07hdDxSICjaKk5M0+Za0xPb5qCMzjqw8K5g458w4ZknFW
auH9Z+2hg9X/93kZE/gy669r3ir0fEoyW82pUdEdNbRFLmVdVwljPRzd3KwLgnC4LGOWWjPBgWWJ
rUqjPErCXFDtIxdxIi/4AGmMhrss0fQcm32dz2JHw54cuzLYEeqzNiqCRBURa4NP/SjiqrX0LpYu
+/tBm8wYb19SEMnkaevVHRm89ewyVmiwVvgyy7Gg5AusJ7gAbXDZbDP+2R6gFL/Quple23dwXMqV
SCKahMyj8si1tY4Ym20ilSsGiqHoUxEcXKY6tRK7buX5Qxh9BDZB39mmYZhxttby05+YxKu61F2q
iiXXjQBbHF4E0TQYl1WpXkHU2mK6nIXGE4/IBKdhLOrLYuGqLGz+/eeGsnF9hGabqSdcAWR9+ilq
jCxHzC/7u1onJouwCBa32kehDZmuVewL1xxRfVTdDpAGhJu04bNJyi5OjC7MJ5hPBj90O8v1vifD
osdg59FbSI5ATXKfvPHW6PZabIXyLthe7GY2PlWtzETpFe33r9XbP0vOVygN6vuhZWQyoiMuZKM2
cubESoBjp98U/KIN4E8ZUlgMqFhRbMcUC8vDMSFvb/HdhG2r+BT0ltDhWpys+aWVEWqAl9LY6OIt
C9K/Xt6r+MHZTdCigI3pHkAbAzQeUFBR6unAo7kqt1PXys6b4KiZrfetcL+lhUi54Wl+ISarIZxV
GjC4PDPTnftaGv3w9LbpV8qK7po96wZrjTXpvpk8hLNVsaAbD4NvJqWu+FSkj+0Jl3nmP1T3XLXp
JCSfO5bF8Cg3SXvg7DX5TN/0HQl9HUsfngP9+k2hagiFoOb8SdI8ohnJ2ILZad9ScWrANxH5KTMy
PE5ldM4CHg5qIurEmYiZ2jJNCiUhOLoJRatJDQRHBnjDAx2pGkOkP57iKopUPj5apV0m1ur4hYXg
20OsNpGBgE19e4ybCB+0lP462tcJqTeTzgDPVrPVOBB1x+oiEvo7i154pmQRoAAIXW0JdmXKbflo
wK499dtf7oWHWdfiPCBWoNfSp5kd1HVlLCKIu0che1X7n43UR/iO2gDXLn3G7RLSnleFNoJIt6yJ
e85l5aNM+GbDP8h35XO/cjbimN7yDNkiffBJPBYrYVtSJKtD32QtMjBtQHrR4vaE5O3H022N5rux
PEsgP7uQ8ePiu0SsFIAxt42yMvmK2v6v2J3sdsWzYXW4fgrjx5qxbVCt+LfSVWWfFvL3udEEBId3
wlrGkyIVUkQdlP2dVv6PSobpIE4MuRNF74y2pQRpM5AgeENM4nTdM3RD+sjxRhTPn/WQLAxi27Zq
QjOkT5ffaMCCHPWtJtGwI2NEMNJhVGk0j9EMr4/Cnoer83HNXhuy1W4L08NHhtr1CcNWUivi4uyh
dR1WvWwel4HxhujSPKfOcfCmjf5KF2EUmDSn9ESOzdPw6p/BFRBPUSDGL7qcbfyMEXar6W54L27b
tFCejZF7fxXablqz8ee6OUlquaWfm1dlenEE+ciwyxv7gtPD53MSJp5k+j/wuD0o9aZ1sgAEPKwO
jl9EbEGEkxfD4Mc0Ox1RI//xm/YE97L8WJFB90QFypabbPtZXaVrQWtmSx1x5RVUmQj2vhswZ3la
IiJH4plqZZIm3IEDk/BlBAMn3n1Zyu8HJarMO4lD/4QWZGeJK4oxEEJpbY5RaNX/Fj/PWI/iu3vb
4b1gwHJUPq/ZklAGROp4xkjTCWzxXBTM0TfR+dhZWWhIOAsgFIwOAI6h5vUXBJLbBUT1Yj5nlFF0
FobqFtzOxohKW8EexiCw4XTx+4XA2li2zAlpZodLRWHJFRowUHcA849e3rhGxbw4FoMy7VuoV3B3
cFpN6PA5/ucEVpJMlN8K2Dj4D8flE49s+6bAAW4MtFxd6AdOAIc1L6bJrrgU1LJjQKHcHgmdaNzg
glE8broT36VdibP5noqaqsXVme/gDkp6YydjFI15R1a6Zdk0LhpHTREVoCiEY6wmcg7gxJC3kVKf
SlQBJHsx7BnEZNJOmYhGKhiQTCs6F3pZ2ubSTS1m6DipOqysqBfYUVyF+o+phdQrhu9L0f6BYTHm
xdHbgFWMrpTtReLuQSFA6Fila7XvsYdaPGY2+1gVVFvU6p+T/uftvEZiZgpbnIS+5flhO3R6Dke0
sS1Uz8j4z/VwWFBT5MyUlgtd2A5SR/raWreviVMIO1WA64/Nns7Yhu89f7RBgBMw3CX1E7Xlqi0p
HzZ9Beq161N5nP65YYnWtlbVUSYcPozWm6ZyxKPR96s50yRmrYvlZF6ym/CX4A6Vt5Vz7O/7cQCW
fVlbzbEKE0d7bAJYOfguxs2AsRD/6HsFq8gyNcarQhBWWaw7/UEn5xKXVaeaaacaS7HAXravQF52
oGHqgzD8qI4Ssd1Z2JYBP+7gW9A00g+YupzJtaKkat3oVgzdT/rPTu3vRLVSOmT7KEd+r63gT9Iz
hmlQsmPMhVJDaqiSrUjKRaZKRBqAjWnTs1Kd5buPzkmJ3G99UKdV1Y1MsuxV81KQ0LZV0QBxizGD
32mYygTiyANas5CUy3KCq3VsQq0xhI6wOIymEtxcytRhCO4jnvI2IwJh2MQuCJCPv6mYD4D3U0U3
aSRTdSxgwRZfycIR90Jy+ts3UvCjmyiqw5TX/6QIPgmAlJbchRTcciD4wS9ZS7/tAzOEdsIy9RCd
jgt/7kLWMXc6ybyg/P9NeCThs7l5+EtvwClBIKFb2XEUAg5Tu5ZRlejcAD64LKpT5SNE+2bUTHyl
yiXA+VrqQqN5BqKt2r356cuz00N4ZDGKr1cI31cf1HtScbjF8q0LxnyS2uhj8CvMb2qqexiy2JcG
bTqKR5wJ3knmp2FpwP+GZtocloUW2Y3jVQgmbWhvVESgxDKh2hX2iyrybZDwqd3MQtquEbou0GlI
6dyh5ycgWJlh9JOFCS7IYbw2DsmndjfRf7N/pCYtO7xQZpGaaNMU3Gahpv3NLRBjrf43mCPgcsPC
mC0erdqvcVpuZ7QW989f3AcsA3gGA8P9PHuXbPmNTz4EywB0a/6Ny2vY4YMlkoJtXhMBjIi3YslS
NKOZOVTWgKETPMxpKws+MQJBQ0TFe7AMPG3Ux3txjpAOFYY5LqbdU0NEsQH6jEZTj13G4JI/S0q3
bhnUNgfXw3mKWfB07un+xNZiWHVWssC2dEYL15RF+hTOTUTJniwnPi2/shXnCIlZWHy/xJACaS/V
D6EKvyisodrEJ1/J6XIpNnjLHTxD9nZI0BY8DER3JieIHbznTYQFD6/8JvDA94g8AEGyJOF+krWx
xtZuDyFQRM0/Id2Y4/NobxKxFpjo+A0Yrkac8pVhHQVlVF23So4mHcO9xa5A4em8pTcmPSqAl+vS
JRqRDafZuEdYepC57fwcRkGGEe1nzdOLKSgwOMFRTJtV3Y2GcMMsLTmVMT6GkFVYsYgMG/FMISCW
RF9bcgcbEIGMc9BWa6wvZIILoIu6dxQTDMaVA9Td3QZNgMTbUXwDqTPexPkqnoJ2eXfldnUeVj7C
oWGUkdK9qM9Bv7HJstUSoKu1a/Pzb/xlsiMCqsUyxt2v48umwaprVYcQDtTZy9LhDx5e2Pafw6yS
yrtz8saltavvq7o1R9+vwgbujpjKF3wrgo/arX5lYDAwN6X4CeblTOeSoO8MRvsYywg8grvDT4Bt
PzdVxY/THcI5vKnFrJM6hxFyyUM56H8rmTkUECju1UULVYaZNysA+k8SFW6s4JihZC0JxH+XONRE
aesveRGtV6r90P77b7jQwnyHMj/7tD491OpVrPAWcaAQwvrNzpU5Nm7/ZojtRjzY31YdAwSni+mn
An5Bq5QIacXPHLBAR5w/MWtAHwOjmNWQG0g1l6Oi3foAPkrH4iI01PxDGJO0sdgmfDD1EjxRoYOt
Scpj1llkJFzB+l9F3zejF17QHBcblTI1mM7h6bPouL1hfyd8+dwTxVZwpgOZ6Q3cb6zs92UCPp8v
1dAAzwA7GGTTFyvBCLRYwUMv9WGEZLEdtQgGW/wjkJaJIfeEnd/wKR3RVwhOqo0zaojYzOfPUWYH
hoZWvrvTDwZe1LlOIwyoSx3IMKbi44P3kjPniueszp2d3uuh62nTmljWHV1i+aj7z9q2AfNWVs8s
iLh5CNm9CGQ+IblYHpGCYxL5CVv2S7MdeuiAGfy9ExEV4mMbn6Y/48s5APtjWZm8WZIoEpva8if1
yfHUH5eriUk+G3lwAQiXp1GbC+pTryZfYk57kPhdyxda6U1ITHl7LyjH4RI+E+a57tNm5ZCgQrV4
M9lmMWUg/5d6CGkFYbqjcwxL+H6+8y79VNQthG3VV8/KG6f/DL6bMItHYqPoSkEa5dEMYpYvGPn0
SCTtCOgSCBHWMjU7Z7S9X5UIRHoK86dJvRwIldocoLfxElWFMSH+Sw+JcsSNAdHHr8EXf4ZRFpj4
kREWIwPaHpzKXHzM4IesjnAKe8E61X0Q9gkTkeZJq3W6NvF8+Ps5KzehjbhsPPIfMCO7m7kgxD4w
55UQ5Pemsnp6Kvhxu3g9x1KOAX12Af8U2su6t3b3hdmoa0T3kL9mVwxltZnt+TZPZ9adG8oxSgyA
PIMslB2qVZv432csv1pl8RgChi/LfuMwz2RKrbaQSssTVaOxlxim2DuqOKME+VxLAqds2Lu4wuLZ
ErvKB19xTLSJV000NuaIOmEXuHXnLfK7svTDJOonArjLz1Lax/W+dLtiVy/mCjV1RrwoCh8BRz2N
E3KTQTsH733c52PM22tLN7FWN5f5HhC/FKQqqmk2PIbetqlhcOcfrpRwXCOBANkGxOpFvHS4+B8W
BEmxB3RQlh0zygYw86ps19b//kV1vPI0twGYUmPvZoQ3ZXpcW46wcG1w67fElK7tDs2dIw6t6OIz
9gu6ucMmRYLpPZzyo/35XyQKMtjXmBPRWSEyJFhTCztTwYHLSz9NTQCZB0cDYJWwn4WIc0mLMPJb
Dw5ZCcQCsG5B9co6jg+tqItyfi6u5fwmDYQMX7FjMT3CyIRO1Cfv2292gwRlDL3u429X8NceX4du
f4IVy2U/Q3Gx5tPredkzNIXZRYBbqFKm8Pva15DJxu9UdxmR1zPmLjswEuk5+ldmGPKD53xOvXeJ
0e5ttyA7NxCCd5E0Wqc7HlQiMMAXHIfzPFamM3Q894FQ4J/0qUkYRblu03s2zzgo/nbwppsgpIEp
BEnkMtf3SDLp3alaI9cUOEu+6aTMAjlR0ie9u6lDaCjCN11WjQ18SmZbFGJx3nsnwgy43zTOLEjY
wer8kU8WGjMSNhlGx0/e+G7t8K11dFz91txhHCEJDEJo/ouNO6ayY55+mVYrUlCcJj97G2LEc4OI
gLuw1zyO+tXPId2vi1iRlpWixx1Pk5w9MLIK7WXBANB9G/xBd4qW5FlpKkwTUGCDvyedokpEuqHU
hBO0hEPArMB+GgfEak2r7kQcod8jM8rzyfUtnQHQMbNPBjVWRHbKkVUJ8fVg/xlEu9eJYXH1QtXp
yUY6laQVv8mWIyxwzoouAPaFjhfQNyLiRtw4083P2I1Py7tE027KyzgRxOUvZIR2DbyO+fVm6wOm
KyhHbF9ofl/M+UwFqsTTQNjdwdRvruLNFXxtlkyN6xCOwNAVGR+LvwnEP/AnLQld1qDZz9NyHdgn
Cu/57ZPpUON7Xa8WqXqn1c78qE3CDed/TfeUS0WcwY3e6EZAJyOQBpBCjjSVcATleWWqMulH2hlm
m8zLHyiV/azt8wwPc4aVW+rN9iciEqN5q8MpAKiYlI2sJIlb4yLHwm205P1kTM7gPrTeOY2gJJNL
BwHydkGIxiwvS2X4YAvMkCU5YsReHB44XbYzJXvsM0GIfSvLkVFdJAtpziXZs3W0SSRX261zQzYB
7n71CET4Udp7dso1Bpd3rXTybEqzsbHXj4Jx/AVuppiTpT558fhjd2aPn8YFHtusvXrkrbFjBgKS
1P+6u6JBKCbN25I4rA7uF4CFer5d0me2CZdgvDAHaBThnG6yCINliUW/NCQjjYlZKbUigUyuxrEd
Uq94QYIOjWr1vSQSElB/5F53GoiNeXbxGgZvA9mfPTHEZ3Wkon3EpiQ9JYvOLGUSeUk+NZh4JJD9
IygzeN7BK1+ZkyPsmCxb5JBtrKNxua4/+06bCrbJviJlJ4becboafRo1a6cpWgNmCNaaAREAkngL
+zZOlAGism/Z7V+RPu+EvRHl1iNjYaB/BIh+1Lj7SLNl7Hq8cSvb/B0qsv+Ncq51Rb0PKI/SZdaA
AMuz/2J9qbKRItsO3udov7fEoWDLjA+hEmrEDyDbj1eRegxh77c/gCE84nwIPs41Xux+D3HL5p1V
DuMJjmjqFl1Tju2zcYrTZMf+gMSg3zorOkDIlQU9dNgyPcqFQIDdF6LI6etaWUET8F74Cdz5Gpxx
Ytwy6uuRh8uyA+07XXKsazTSPat6DgxdFmWUs/M3R8aDy4542gD5tRiG1hSS+pwacAF91xSccsSi
wc6LfifVQehZ9T0PXsdkREx4tBqDNNjdhXi3gtb84Q9OIAq3bmc8W0M66UAFaCivFvb2lSWpWXIL
e+ZAmRKxJ5MOVdk9oWQDRtZ/ySeMd/lGAyWaQ6h7UEEKoqNOO1//UOuMgJenCO8QmrZCnVTJGAaV
Gx2xQ6zsft98mYAsWJ+Evemij8GQx2j27EOvsj172DJ9TM1nNs6DrSSs6AE0UlfAfd5oSjYxZbQ6
9BcyzNpwS23JDhqH6lAjV2Dd96vxETPjH63B0qLhLwVxBZRDMWuYr/S7xGA3VT5sh8UkX+XEun+T
yKONg87F+SZ4DsvtBeLmbiWUEY7o8tc9LKoKI5rIAtlG118AMz54z4zQVx502UJjZYyDebT/K5L4
eRU2ZeD3l+TxquyAI5tYfAmX29RID/vS4NUrFNTxEAeYsIG9OVpIYbQ/tNK6dFAY/h13x8vqGwkZ
HmInFhNY81q0aI+o+IeXP6sF64bZpV3oP1qghvofON751CJgspxw3dptJcAFmwwrissDN6mvURpV
RlUFYdJULpjiD70RiIP0cacFCk3Oi6W58HOkqjhKykwW+y+W1yq1o0vH8ILRiLgdA+q055w+KsRa
LWS6ah7csrlpJd2ioey+gBlcyh28z9/FcrhemwcPVuBtA7GaNu62mqfW2Err5l7qxJxepCDXY4Sa
YUsgaWkcn/JKSHEc8yNfgnmWcdzIsujFFq3p7OiH30rwqh0vjaARAqTYe/Uum5Hy9EU+Ay1jm9nE
EHoulWELoSCyB8pWxAr62fw/x2kbWQkFMMhJ/c49/FRp9vFywTh/9wjfdHXMv6/ieOwVKpdidSYm
pukxfvvZfIXJOPAuYeM5lpE2L/eYiqspIPDMvjasLOOkSW80HMVESztwCkwAbAasiRP64xO0oCGj
e8IljhXx/Yokf7ntrd8+uRxeenNzIB2Yx5oGu8G/bQHs3Rr9EEQi6bH2wisccBAxF05yUi/ieHQJ
jELJfo9zqFCLqNwU9bLnT8/7obfFeCaPHwrykjrlXC1TksLH48lhKNIBmca1SKVNjFtEYMIqevgT
RE8Cie0VXTxgGH0j+pOpNGL6PgQ6BxAzbbXc065zAsrbSj2nIP9520g901QQBmfAejy++6Cw/Lod
/QRRGxYufuzoeYk7zOojWlaOQwz15RHyelyLTJT7oPn7pABiBhnpM7tKIf3s8JusCnkage3J9HtE
pIx4GBXKmtgl9Gb717iaQdwFUhPOp6kHBz3oZ/it/dqP0tJxCcNFZMZc2FrbTN6UdmOASqQA8R+h
zxpoeSkp1GUZzpO+wMGgPiIVxs71rfQMW/0njvpjyo2uEMHoPQFJtbjCJuIJaTBvGK7dAey/w+zH
a9uYFSY4pX27/7WbFZdZfhwNWIQ2tOC0X9xWB5xpOwNaPu/cktwSevq8BN+AxTIZZLYvVUnFYqSi
KQc6LpL133/hIHYGcSvv5z5l9GdcBYM+b18eNabln6P6ruy0YrHVla1YKnatOVOIlH+rbP1onfft
C3Wu06eMF0MDbnIdLASgx+TZDPQqZRaLZFM4ATeSC7yTB4dhlZs1cOCN9zvF/eHBg5PeQHzdVjWT
QLbvI/JRXz+0ZVFAwoomDvUq6kx20itIStELhFDfJywTueg+RiJFbsDpCpQPVtd8K4yu+oFjfin0
I5tiv897MVS1cWU+BIuFYCuLoI6D9CjJEOJDWjNjl5Fo4mXgLtGaDijHguoo/sIzSFU5Nt+vA/bP
VBPqwG0rt7Mcx2ftfhobb9wlQWjnKQ3+rIAC2v0WLhDkaOeFB2xQgRTa6SmMYOUmt86jjFhAzkgf
IIjfLz1lRSyTdNbpA2kPaKifBRq4JyJJJTOpzRN+Fhr3pX9zdu2Wkkg8MYcK4XtO32xXamRvVQAC
TlRcSo3uC14pz9fPnaEZFWP2OmJ5z5Sn8W+AyVzPxHTdpxfVRQrPljjr8xrPXJGCNK5Ukg4V1pMK
B8B+Tnpe1F5Pex/HQnC3qQXDia12G/j75HZmvvxfPRuN9ljei0KGW/+1lznqyY/ICg4m2sdeNOhF
DC90Pz5n57mV77HKMzxvwQcZ6sd2CHrGitIiDlC816iCZ5jsep+aJ3IuJOtuFcQKbc0FEUuoaQXT
R2D17dPjdfxrxE9u6gikemofTujau06MTSXvOOupILXIy5Tiusd/XOaAAu6Jn7GJ0b2dG/b9FwOH
yQLP66DOtOh5Cl8uFWyY64TLH7BF0kyxmzwJxegkg5lYmewQNs1900PA+51V73WbXOmwXXxh/9ko
ylFMRV8FO+4Q12q/3IFFydSPPcvcDdBsbrjxHIqn40tOs20qHlibSdqsHXpvIG+CpRnxMyyxbeKN
k7E5dmovoh0LR2fZybbX05bZdoLrsT8/vOZHXD380c8m5BKq0GMxmj2hjKcmdl29LIWAP/Q6I5pk
djOX3h89lIBpuU7QO1TCBlElT4xYyvC+fjH57FNPx/KQYATS5XfAbMG8sOL5sDyhS+s983kyT48Q
w+WNJ4AYpmVgdndFMPk2GlKNPtED3ubHsX/bIMxEtNbpEc4+ModaUmW3kf3Gcltlh/ct0IIwBdp9
Q5UD45xZqRwLYooi6o8P09Tbu/fvfLpUPVBvp9KNPJ2Rcb+Sj+a0PIaPp17jrWVTCZDCX/4lJJmu
QEcohhIFkjyf8idmRBu3hl4p9lD+bi8wjek7BX4UQYiVz2zsxmX9wMOiWvggHEbWZCC2xjyuRduV
SnvkC/11lGA9xFg/OjXYRe9Mavr7fGpOWdQbBIVmEjmVgpOJxrUu4iB9Ij9yBh/HP/n209/1ENTH
JYUS45n4Iwy1/jbNKewGDGjwYe5beEfjqA0DOHqUCGC519tzDKRSfFXpomJFAvYpUD1BRvarPcbO
mjXfxnDLydcrAGS7L9INNILCVaaZj5/KTKAW6P18BtC7kBXQP2ZoH37gicdOWrXbu5xsnPsjp3jc
19j5sv0iKPWcnKJMjkXrfpNIjvd4lI199gmtz8Y0Gns2zwKIr5eH/dQsQfYe1DxxlxVXeyuVQ0qn
zopj3jfi/hSBQkS1G1Q06CpJQB22VQo7b9U8Bv48NRq4juLSPeZpPsHC+NH5uj3s9WhYkbFN4dtu
hhlar3bdc726bLhRUmV7+opULwThYl3eaP09YeYnJXD3qrb7eCW8h0rtlhiPvzqC2Y1pg3dTHsX8
1Kj0TkW8JNYp78+50FuscxGCoQFS8C4yS33PFWFZTBSNHDdeGmAzyTsGBfxDBzy/6lIdHXx6XwJY
t7nacYwVBwq5X8TlIqT8UWsli5ObqqTak9oAvMK/5ZjkNLqExFL1/motFz4NZrEVpPLOGOozcLkM
QsWWC+PjpImc1WnBHxF0gQQ06nIhJH13uYbfJkMWh+0EZ3cwLIoT3BCxYndnLwzBv8/FAdnhJNIj
CfKHRvUbi46gWvo80KqnfJl+VpqIYZFc9t5Ri7vwYANG3G9DRJ4P4AWtGj34bqim3+b5A5SPY0JN
/t5LdUqPHJo1zMzAjD3Gqx8ZSwgd5QPjoudxmj1/a/iIPopgC4ONTHuYaMS1NmyNFEXFbOWzv+Fm
Zgn30zO1h16qUoTBHb3tKTjNd5euUcz1MCXiVEY/jpl8UDD6dxQBS9Bf/lh4gzblE/OqzpzDGifD
7QzS7K7vtiBavHSj8RsMue1662GgimAJ8esH6rPQlvJFEwRyOPMLHXsoZ8DDMVo8UbruFelsJz9u
GLZsLRocD14Z/aQ348ZGmolGMJMKjltYZNHBewkJ7xrOC0t8Uhhk1XVVIAR4S9UhHE1zW9mGRZTv
lB8XnyW3m/xGfTcqEERtnClfOfI13hUpGCbDj8xKEDxlUU+KMrmNx+E+Njj3D3VDLIGz1DvM+8+t
q5LOVrwFhUIWKMq1ybL7Y0PiE3DPZJwO3GEYSEVnWVRsEcunPEfJt4Nw8rgU6r2EjZXOWW3MZLXv
CZnX7kFz9ogrlfn4nsZgih2gHaEfrjs0NYPYFQW3aGa+6ZuV1Z6CtbPn9X8cVCqEpeoPSv+LENNb
U0kjLMD/cCaXolVR+3AbsvzxNyy4Pf72iKFdejPkBtTtYolUhSzCpBtGGpLURJtP7y9WiCGbtRwz
rc93l3cK6gN9/0moYAH5wNklgKCB+/EFRb2uTdDkpzutAm6dkqY3wNM5Dwr2ETrF2TZbce3U1GRY
0C15o8eID1Xx4qeD/j88L+Pz1qToTNKMzFsMHrAlxQRksyeFdVdsw2/t3BiA3KCM0MoRREZZufeH
pnKQUrY9kqfhk88zBkoQdr3yc2GdTdTIkslDXHxQghGqkrc6YCD69LdljrKOOCKUiTdqG8+buOB0
ubtMb7OtL8WIJ4XDUzTAwsQb5HQG+KEvHy2LZSjBH4fMnvfjC9sXFrc+q+bQ47T2BrhO4WY7OWlL
WWJCK/9aEvhHTMwN4uKuFigOs5/TmjihB83uAd+BwpScZ1VQzY6OpKhM3NQ74lxSghHqd/f/3oNK
XgC90zTIBNGexG3g5aJzqLdGQbbQCySm/je3BNajlCnPPWb3MuAgnAk25oQFxV4W8lx8mBxMYmxe
tXpMRm/oE8RfCIXnPcc0XE5NoI5CVO2T/OuaHn9VRQepap1NYq7GBaMTMoxddkbl2TPJ5jEQNOyY
GBBwnWQRPbTESnMqwCjgCEDi3VdR92Uz3tTedFndkG4eeL8dVuj+h2y3p/4tjt0Wm1unDfBBTSNZ
OdN8c4qEHB07u94TrpE++z+Of9Ih3Ntc0V6FB6Scgcud6HDqkgSuY57AkaagNz9KZU4yV68uYlpd
84AZF39ZNcIkV6sunySLEE5oxM6uWzm2cq2Eq+Ut0oGSr4s+M5q9hD1ooTehONpVg5G6Kd7v9ZvF
a9HDLDKpaY038FKuTO/2z2KoI0mbv4g5AOjcyB9dsjCpAIuMiRfdbElP8EoRMgp/ZugpiUquuVgg
maXVXJlgkmP9phIEGk6zRci4OM+IXOOqMjlWSZN/WnydATdCHuzhTcQt0n6SknBEws+6gOWpXm+J
DCP+FN0JZ6rn7SvFUMVnvDa1/Vlz3CvHe1eRX8J6ROZ2gvX309ELMBEbJNU72BJ50XREtCIiJxPO
zai6V42KstcKRLwfsDkARGBjMv0Rb7Ae01dJleMGweS/9Zo41MShF1HUriQ55e4yergUk8h1Yru1
ANBerwf/v0fo/c3z17SC3+BZ44m5NvH/fK8vzsbuoZishAQHuZ66MjrxcqobHqWLcpRVOg4Gejcb
TT/giAZ+i87laDSY+Ugtp0xXRP2qPaPmZ8mYdv89eg53qxclxgB7Ztr2y86g11F8L0YGzhvLgxHw
PGr0BQDroNsSW/QaG2S+TOnAzAV1SBNrtVlf89L8gKdnGIK2GQLIbyv3pDzNJ2+G0KHyR2zcf+wB
8CESyx+MDnIiTUKde1nbOEaAidKRhfiHllzil1we6FNayVefSSczLUZ6NXRbzOoT7Usg0GDQbfdM
UWd/OJaA1QaWd6x8fYPs3oGkqYjizOPfzU1FFnSNj0k10pw0bF+apaZAt1aC5dn8O6bUQw2tgDDa
rIZGg3vjHGl7a5ZtkyUPb5/YeRuJ6I+UT+dBGajr3YQvFoQb7n0pnJjfdOE2f0QX1g2FHnuZ7x/8
xhYR7pWDWRhNn7sjj/xWY9mKCE+G9g+Qru+AewkhEGCQ+18H1OMS380Geb11lpwrriSa6lTC4hQQ
994ET37G8kKkwBuGyo7rpb4TNYkYHo0RpB1V1+bVXU9Qqc2ZlUFyqfDqjv5zrRNRQaxYjI6kB3zm
WtKrqrk34XDLRa2JE9z3/6/c4zzdL3W8l52bSV/eTk+G6p2QbT5oeTifqb43uiDCyUNiBvtBULjV
nv9McMqLuycwOtdmAc9kzrnW5mhbe3Dqs5637N2x0doM0SaNpE4U1p3nXozm2EkIoYtIpQVjSDVr
cJ4P6ZOAqs/7Z8kv6QAPkkxeqiNl9TnaEIGdGbRU6zQBi4m1jK/TBEyl4uKL2ZiWZTPx38s2G+nM
dfp5VxZhOyice1oKJkB5+3S7ytajezWsX1OZJdgjW4XHeysX7OEf0eiGyJoYOu18Enxf1Ka+9JfL
uATS+nrasHjaMCdt+QPxTXrP2CqhuK9PbSb1B8UAOy9Jp8+hzv+bmuUjqjkzrIlcz6oSsfLPskdb
+d1AlrO2qUIxF8kEZyiTWh06hB1sgpP9YwU9/duP/hqiRPFv6tv9AYaFcbEHQuvvxPKzkokRtohT
DSlY8CKp/syksu1HWTK9HamkX2ZJ4IK8Y0xVN2VKdwbUXJIHLH0TaZ96GORlAjyq42GlKnIjhMlr
RjpNYOqc80FM6FJg4ufvNFmL1RMwlGlsEF2DYeQtzHdNqqlgUuPcXoRI/1rJjaoC90/qP5thjh7F
f5aCvuhZMpOLNni2oiVPcHQNcJ1jWk/HLGKBLmo9MdspehmNQ50DBl3rwWHx+3ziZG8/Bh4F5Em2
uKJlU9WFyPu78Da2+EDIi9HrB892krhtFVbYAxSk5Vklrd8BgyQF5Amrvm96JnuQ1JejV6T2ulLN
8HKdLYcNlRwAG/ebr2wMT3PQlv6AWs7LLNd3fETfIYPgu0eDc4QSbg2fPV84xczF2Pu+92pynghV
GiNBzOrFyrrajDdpzt2MgrVA61SKTnsvLiAvM7AJ2rfbN0paXBUkAK/DA3UJqK8x1rm8ntne9nYu
BCmSVZEvWwl8elmlc22lTVBrwp9S96Llgc8/aJ+BCwA9fjw8N2Vrub/oRd76U+Tqi9CIfa2oRbQ5
kdkoPpNWp+5iCt+1GigkyWi0eU/1y9lxStcgHJPvXjzz+yoziyHBCAsFBycOmfVgWyOrg1pULKPI
KZlBXwRUyJPvTQ2URGJRwo34KVPdGBsHm+z3wlFpkw1klSkl3zWWbx5dL+Wy0eQZMnoKxxGOs9+O
NYlVP+onSaZAwUK7GeCgzq61QkPJ4siP9VAuYeAPvJF3CJdxB2AdLwhRQHCkIzE1r9LSmCPgXerQ
UqyKbtuy4hncBZ8JXGzLSbRxOPEmFU3xK2HRsmWiXtFWSAK6+LyiBEWATkiIWelQu8rnVPYWNnKP
bcu5MKBGYTvTzIIPKwV360V4yY0YBW6k9yB95GouzVgmLEJlgPcCgsOlXq48j2rKp94rIUZv+ojG
Qb/G8YwDUoFwqsLLW35hzTYxegnG/BlOJiXzf5Cqdwei69oygP3orR8dhGDrhy7vFOtbAFeJWZu+
koXmCx/6HE6fIEiKWfgL5gjZG3ZROL9ecYNni+vV+cJVkc6hIPTS4/YnG6jBjpKEBtVVLEv96aa6
Lzq+BAO/dqFexy8fh7uB+D8yTRzCl2hHIzcSyxPKVk5hSBcKYe+bW/GT67/2W5skcr5ayivxr7iB
VErBPB22LF8n3whP/1BNbS4MlhW1VvxXYei6vRDWNTHothv15R/JL8Q5ckadG7TLLq2iICbMU33M
4SOOHEyMk0Z69/vKtzgvhljQqy2BciusGKA0n3ru7CurwavvRWztjlHYliACqEkm2b3Bwkp3uF27
jsQhNmi7mT1gAfNleJtD2ceQLzT/nySkqJDZQeK61R/WoA9P2+VfunqaVhnOBECV3GLxcPunEi7Z
CTgPnvgQJJ7s4nMqUFDuYO8wWT1s9nnnEP+eq/ekEleBtzZum0xu6Mynr9KpIy7j7L/TPIZRUBLJ
ZVyTNwQ7O0sdEBmVJlvgkpSQsJULCmhNj62FPhcIi76ca4s8eq863VB2R1kFaC/EaL5w4IMyPrQA
mk9a9bCYWA7W2gLPrdAqyZtzYYPNpHmH/6wXKAJI6fKR7kavyS/cjTqr5RkJX7CUPCsJ7nP9dW6R
WbSAMz6gar+r1mp4I6v4jDWQd6JQfHiEGcOJRRmO1N5Yd2UNLobpP6Gl0xLCTQCtXdIaYIBi8EkC
rmH6+sV3aQQsJQrXw8W+dS0nBn/zNhd/X+cchwLSo7+3rXFFGc6TKBXwyWwYHP8tXCRZmydpRgGf
6splMVX2mDGtfsQjyXBKB+qN9qcbLBrZvRE3LdAYBE2bCeU9XhbGmwB+JMsrTFvx/x/oP/xus1bE
7geeaEBS1bREr+d3tjSdlMLjN65XKdDIci4Jm6RZ9tAG+/fX4wT0ODNfe5cz0htNszamyena+3On
fMm7VPV7j0bJVxysc66p0SbxUuq6jNmO5v/1W8aJnvFUHsFY0CYxnm3YqNOE9BwQ4R9P4qbQqFLs
bfzLNHSxOEd879LCKtKtw5gr6/2krR0zUXzeaW14k6/eQiA4rV9Bx92z1DYzXsHbbwFzO/Pu4E/l
hQJ1MraGSNnhjGDOkSIiNQ4RnJ7HgNnaDp4wpWVl3SJ5YFvL/4CpYE7ZksTyg8/OW0kbCe5/yvKi
7RmqtmnVURlM05gyF98lm73zD3ivZf+VKQzA0KgmGyUTv3Q7EsZoMPmtFHpHQiWAQNc+f6fw4qm7
e6fRuP4i44L3wcacuESRW9YOiRj96D0GrcNP+hKewAZduNvScEHCN/jRv4/YiykZbuxhe2CKPzyM
vW7xMR383XPR263H3VTrlMMNF2AANULcBix+eWXEQ4zGaF3XuURTr9jD6M+ujrfsShSI1L6228T/
KXan1vKppqMHW8CmwYmpiWKiT3wBVyiomkPCG1feNdkB96KlhiOUXnAKqueoeGEjOLFKfIrK0Izr
ov7f0CskgfJkiPgl2tv+bwprF0aCOK68DZ4xglvln6PzaeMb//8272BBzIaZoK3X3tbtlDzSHL2W
wPaoooXU3f/Zsnwvz9C++sAI9DryIQRATcFRSMKKIWFBP7m0vNuRoTTHCOa1MMjlfT8yAaRkZh+R
7DiYfkB6wePSbhcf515AdJC50ErZ/Dz+LpxgGWNrxzOHrWhXQJSv/P8asYw0vf14uoAWV0Sjj/vT
KuoGa0gNdrPbIUM8IwVTPpaKYjiGwdlncJ0vBKfc3nrz7DCA1VYQeM1FJJrAlEr0NBzBW+xXlyLq
PfQ3LV0zSEmECN/vqSyQrHL8ZKgLccqt4NllcV7U1GTBtredH7d9j1babHXXtyBt/jBP7MP9aA9k
NVQ7UOJ9xNPm0JakzKv3Hcek/nhXTuhoodRY6ban5SiHQVDa4CVILexe5+OdgZqXqdqG7t8yQ8XP
B5Zzv3idV0C68/RQMEf5+D+693tYbse/2U6/zXDAn1g9P2PCsom8a5Duod1afu9ijFcfI6IXf5Ax
CeQHWmCarE9FR9ZjdigY54zNfDXHy/nbIV/tGhWVNrb7I6PNu0t9g+rpIHqzz+PyLRlznzJ6Rbqo
R73yXPJJ3/dHHbsQVA9qKf5cvOy9K5m4tU5s3kR2Sy5/8Nc2qRzdYFK8fuDNEVThRVqd0DwffGAV
37L2aliBFtqZGqYACeYCZEc8tVP3gjRNnS/1RnO4qjnMh9M+woseKtXwkEYYtrPg0UfmsXBmc8hX
m5oxxnmNtYL3aOZQL15KjcD7OCSL4cghcdcpaqjd+uldUNQkT2KBdjvvkQj1uzJb6WyFFZJAZMji
n6zd2rygvN/i/5MNlWYgDLBpfAmvlNw517reultJeYT9ZPKigORGRqis9gj2OHfhcWxOZljiKuHr
PF9G0WIWI43fvu9uZKA2CiI06OrNRFP1GFBrCn3yZiRSniQwfx/XHh5cwRB9zi6T8HuSMke/donK
nUnmmZYGgGrlK1pEnmYJafDC3U9WnsKh5adVR+JJWQivDrtkk000tICnd7idmXxmZBauV3ZXhvet
RZ2FiUE2qTRHHn3DkwcGqE6T658ED9ZoWtvOilE/QSgrdRQ9/5GTROF+zp+2jZRB3+oVP1scIR4X
PgYWqfXet4zBeisS3dFoxM1obeA7YEncFYGfyhC3496u3POdehkF0Sb7rBThiZzcsr8NbnOlMRyH
DIwhS0cdYC4hveXwcJmUPQsnNiEbouE6bmd7/MmuXWq4c8eZM9eHwl52Cw0//mbMUNNi372gq1/o
EDd8z+1Z0DdauzVukI924f46CMgrm6BZjeyH9aa/vnNqInLQ5BcDIIYqRfEt/L4WeMNKKwfjm2jq
qtErgCyfXXFoD0y9EynEue1idjB1PRafBXCFPjpsoVP2rKFHjMvfieUFW2l/s2QWhKrznF7wYgKI
tY9in16JLUqMnsnzukPrVBfMLuF3omswNQ3V8NfE1RXQSYK8Cibprxzk9FtAYgKHAA7EUnpuAf6c
3LQY+Q41ZGe/Ki58/R7stmf4sUK09OBEtLofpaBubgd/eRb/1AHi1UHULF+vYn1NZJBsCDna5jD6
sSh+4LRYtLJV7M3CYO/yc231+qu4qCIP+edCNTIsgnOhUx7o3RoPQzF8fDN6Gpw1tWms6EZ7VEvR
rF9fTG2YNkrEn6hdWPMy95P0wg+1fcXq9Dx/WwmGhZThElXlDwasBTPVOj7stxTeqETKXW3ftHH7
TyIA8W7mqYFEV7Hn44XYanBHqIdGEDCdJtikX1prCC6dZhy5A5Qd0svESXfn/LcKYUiiLtHz1BgP
zaGoFwmocMV1uxEQXsKS4rkjOOFRD4RHaEcNylnD1p5wyZg1cWooVJsndhRO1isujwWkOYSEi7O3
FjQnM1wbftz7YOLJoa53kL0iXTKyyTp7oK5MmpnNm4HMYR1KoVSfwM6fDkTeuAspmoUxMrjIxlyl
PGoJkM9SnGi5XLWZ36FtWTAEDd/ebDW/dYxu3BPPmE5BfIBYgNJGa1D8M3frFY7r/yoUIIHvKtiK
a9LZYvc/gSlMQzdjkq4VueqfzMqnvt7UNc1y/R9YPMRrsh3BSqgT1VV3Lip8YwDSWqJxXEZBwWYp
TKZGprSXG7qi3aoxrfiGfBOzEtawgD7QHy9tIMd1oo3RFnnDcE2r+sDRkKZYyNu2oWgSu2oSJsdH
aM5tDCHOpvUY8tLIlYUlEnYpehmgACaUyhP76PpSJGFs0qkoQAuqp9GePl6sLFXL+cqAsCVxpkLb
sTDCVlxCUFSemm/z9369tlc/sxu/K1lQoqkAa+gJiC2Hl0nU+KFyse2rgPOwT4NwK3Q/Wbq1m95h
3YEyItfnYGMO6d5wSUrBe0tlqdK4HmL/hxAMTqxBRc7vyTqocNsEkvt37o8z/DshJkjFwYs6Tgp7
6ITWIVQcVV+4bUBFeT+FN+cFv7+irqQ5O+bRlhWoTJ32m4cRkNfIAt7bmkiMNwArwmEGGdAx98HQ
GZxLMFHLQj3ENRZnM44kQE0YHVHpEyjJGJo/ihVYY1sSub/zvGxmJFHOObfbLOkcpxf52MtbX+fi
l9l4vqtQlIDa4c+NEh1HyLsVbKAueJhKM98YfLbahy6XmzqYe25gDZD3xdIQoTjdoUUu+2FHGfs5
Azmc2WIqsaQhugLwDHOJ8dr64GNNE+ZBnbpmebAETp5iDcaIrLd5FH4rE6hUAloz+kvaneWlmJv7
CqCOBfjwxsATso1CyJ3be3/MWp/mR4/l0oB2KjVQZNkJOWW26Ee4M53ALi7jL3Pikfz1feqdzkB9
qNwnwVzVnD6pPGQRh26+a0qoCt+p8Rd6gt4a+JWJ6vDSNVsAvzWufyLiZu+/wGywL1pQabporOGI
cQFd2tPPxUBZKW117KqOXaXn2oexuOPlbbJiRR7ErcApMRpraXptRxw+xmMKJzA2k8J4Cr0+URtk
zVDN6jE+VeNmBt5NrBeut/JcL0RJEuHphoqmvuFce+1GXPGIcKkRqlIAKyrA9jULD3WKZMzyL31t
RnZPv+YRCebVeDgp1l2vXkl5F4RYgFo+GY5NHVyP9wbHwMZKz2pEpFfovlA/Vxtn/qn1o1Dr9zjo
wR1bziTZsTsLOLYVINE45eGH7+G69eRcNBahVsO7ZMlhJjreRiTmBmHVXrFHVJh/bX5qrUFOOZLp
swkDlZYSuN9LBJUuZ9VYFE6dmy16Dyj6j5ac0qKA01hqYBiSpnLlvL2vb+SlMF3yCCWKPlj7RuGd
jFduZKsiKjZh6eU13dx+Zs6ncHTI9aORw5Owqbu+KQ5r1hFnKnmCp+/MbGD7EzpU0jvciFJMOWJH
7/Oc3Jb1DjCRbesgcE6doIka9AN7oi2VoDUY5fIDQ5W0XPwLJwt+2imxQVX5H4kmDeETSwl0kTsH
an9khIHXeZGDlP4tnjgtgr2zUdq5dv5+QObQUTyy68U8p4yMkgXudHtnpUQOvP9XRU/+l1oYZ7J9
XOsQG4x/pkXAOfKodLZRghULJ2iT7OSBwqu0ol8kw8EuAdY7cCrzYl3d7QF1Jm5rrv2YQyXgxFCu
Giespg6QlCkPEefboLHntDhEPbm1jxC0RN7CoU2aZ+ez1zEFu6h79IqKwQ3sJunvERPMBNb5js3A
hm2IARxwwH5mwdCeLAVdcKMDBT+E2YJjZtMCsiQm9YUJswF441vf3HFvlUksMTMjutvp0siAWefW
kci22S07s8zqajxx4zC28nTs0x6KVkgb12s083p0VSu5vG3CM1KCmXe5g6CV1PHgY2zOhsfFF4bU
eDKRenEd6v8JpKvQidixTiSHRSce1kdUyG+I0dxaoIQXI4HPzjKQ1vOqagxwK5UxUbb9X29dNeCa
cVrK0FPtu688D4GKui4fRuiY2LOo8TLuy2tSKXanMCnz5JEw++n5FfRytk4ReUh/vSK8bHliaS6I
YxCYwdv9OLTEsqnaZ29iRT0qvfpgOmV2Qo07TcocR3rnKXfh5R/ZKnL5IebkALJCOUvAfSdz0BQq
tBb1eywq6L73No9/UbaZ2W/uC8PWl9ktUmAoI7SgR3WbDbrEYEyOONnxMoK7+IqoAYX+HGMYrP+c
fhOonvU/cYt0d60dUl4xo5RvjkPwSf5LYY2dt7pmBhtMorFRhN1stLWpUreBIOO/G3KgFTn7gZO5
AgPttAhwvzVum/fpSryLHaCmLjhCq47yvHkQr9UXzKiIHoqyGyQsLtz7cLu9vTcf+VAA4ChSex34
Ma78xgGrxNBYV14hYHoQjnZ21zZKKuYZf/xGZoscwmU5hHmbXjuswJDkyEmZ1yzmJa5Y6EJSVL7i
dYB2u5zIK13levEqIs8yO171gSJboXUHhG8GaJyL72IVtpedqKqmFibzzFFbCh2TPM+120PibBoZ
+k3JywB0JVTRBTvi9uSuZHJQ9fbq+g19Qjtus2cQXTmNCZZL0v3a8l8ttCqzceQFQ92LhH6IwUIu
nDdGquLj/elsU41EaQomHg/rQXla3foZ1zLaBGoy5YBZbghOxGARi3jFWCLUjUyYQA/pp6pIpriR
BoDD636tN1Qh49B38wsv8QFE/apN3WpqnaBfQL0f0kFQFg0Axxv77Ges661wzNSWv9kHZI8UIMI7
8ZTa0I2v7ZKgeYAUoabIcJsDdL6S0gnOADcUMiqTDK+nQZU0I0Ue83u3kurPlKy/Nv2pEJsqJ6go
NIipTrceB4vGxlgW1ysZ9F+Yi+89rcS7Ifvvf0yt9kFTOy4+V20gHqEwQpzslDF15HPZkgIB8K/e
Bm0OSZ2PO/FXeVM5adZYSV+h4PrWWQnnKu2WVYQig4+qVGo/Up3eNMZT5fmTk1AiJFXrx550iE2H
k1lGiOYbukNG13BKx9vInKVW/1lnORg/K04AnhTOHzW1lIRxMxSQjz4c6oUCy5j/aKtXFpHOKeeI
7EWOnoDZOBwJKKUTa6sXUgcwZc24/fUEOTT5Z56y1SjWdc9MXtTbnrh6pt9G8eJsLBtAKkDQW9Nd
59F3HvyqFReFjQQT4OGl3SnNsUuE5z4OEniF7z6lXpmP2AG4ZI3ABclnmtx9mD31oZWUiyXsxeBe
IxFc08XWRC5mR6X1f/2K6LVeQlPUFADsG/vs97FSfZVI5VZvW0VLLy5wUO2HyKK3I2wBs04I2fTa
2E4TLqU1sUvOE2x8boHG9bpRJI2eGS9NhIBPaclVjlWotPsdqx9HvqsrJpnWcGSi5cjoFIOxJUjD
oLGe0MJuBu14/LSmsrya2TqyEdNpdZFQPC42hCEjHHJOY0cFN/4DnzzsJ42dHdMuIDbGtQvsh1k6
7YeRhtu5LJF7f+Bu+pEgZ000t2DOs3pgvSINeftOFH60E6hoWr4LFgPOc1sPD82QBzu1PK43nosf
tGFYG8gNwDXmhmQPH+XQC9PdATDf+SmASPkw1wHG/ojZjTaSpYKf80FZO7JPH1tReuDce2KfOcki
phToR8mweeB9EX55vvtzZrW7Y/bs/fMjAAl/D5IM4fVYlSArZd8hNuHFc23OGLqRjKKW64peP4UY
KtXQA9DIHCAeVI6E3OFUFvBroHOSU1VXOYu+6z+sKZuzE1QeQQr7942QAcGAki/ORMMKIs0RUDSL
SVkXBDXd+wus/M9lig5b4zDF9gV06Ze6Rd2wKxg3kBpHNUVXKaicpD8JdspO2kM517ygRYeW4JnJ
7Qi8wqfhNWhnHQhCogwIdsykQWizhhw8GZZCA9Qaia9dfnISXkOMCW/ZTGAi/xL1E2Cozc8G0/IV
Y8WpqWFJCDNHQZg2v/IzEGfrfZyXFlU/3lpNBEFlSHWdVLqV26no/iYl+YqGHdt53hZNUfhHCKSd
DJf37DtlN+KUkPp9ldHyq5HJSaPexoqPWeHNvHaNfnbtMtOJk8Qc+nou7UYYqik2K6XyI9zaJoKC
B/Dq5gae7ZWitteRBI0Pt41rDdQbZhhPpVTlRzfy1u0v6gAgQ85IXoCPB4Nj2Cf8H4GEnbqj4HAv
557hfsThLt8C/ebxQGiJQRcevGeNxjjeqDyEmegKy6knPzyB90hMwH4lf8/a2j1Ce7Z0ncCTiBWd
UtklXvNfXyn423PxCPHzgD4MNQwNBye3vxlR2gsNvLT0pHOLN2CbctnxEADkMedCEZqs1JyhZjjc
o2eebd0KCVqBhoCfuiKYbm/V7Z9aLV7iODvKT50G1V/0emG1iczLqX8asHV3ZLoJ9GJqiTSqTIig
SK17YTBCMyP5vht3yF+hDhXLfEo2xqw6h8jT82FmEzFAyZumiMcEyfdfVeVp58KsznWregYP00JO
Mxp2qluKrPgZoxwpbUedqGCv7rxQnmNdJD1v8FRkgtjTdM3cFffnIdBz4m2PkUd56jaiAVK97qQ8
hhJgMQG/vaH0h7WzjQzUCmIK+cE50LKdkttzx2VcDEqZZkgUDB7CimskJDU9Fgd7IEqJWMkuNw0k
alWbng4BkhEkRQNq5st40xumz8OF0fQzwqvJ7x5LDJIQWV1sBWqN/JU3d36TIgqu3fvfUJnv0bK4
+mRFzBjRkCm0I8tMMxCoi7knh0+ugZWi9P6mYaacbe+shsu51qblUBLUHRrfwxXCYX/ymb3TlvoV
L6t5ZxPNwjhRYD89MO8D83YYrUxTp03etT90As68wKn1ONjc2cPM3z6B550ph5Na9zcXH6qCfjJ7
BCTJBrfTZohjXGUppmh3Ek2dVRLgxwTMyD1u9yV11HXkUvvb1tlOnI3+KhHAatVEhtAQPJyybsaP
uetgNGETXsafEfvU/EdHuYv8GpURrAeTM2xgW92REeQI5f+FVxNV+N7VUKeiArZhHqsJlfRtIlRo
a9EuQsQGa3FQYoJkUFp5GYzJnOVPamTZpMu2olsIoo+dLvyp7Vl0ZTEaIi05frp5FTUgwGQXlBc7
LtY23y90k1Phc554IjNiy5QOXMFcnzqxS06rGaXvFfGqnduUZH3/mnzqvD3A01YfoFA9roUhG8VE
cdRl2MLN9oiRPr408x3EcCUQ9rHiqeV6COxQw0qsLbpjgnuKfUe4NbEKlnWxWjqq3/gMo/7Btv5i
yQyBVolaqTiN/ttEDmGRYmNGvyX9nxkscE5AIBsREci6K7U+l1ktDAaUQ4knBQtSWozuIW2eBYSy
E03a0XNAVRqbnFkiE5zULTiqrEZCSScKf1mhb0RSFg2aN8LbieYiVLyR7uBt+n3ZuYG8kNsXcQHW
FvInzP2iHTXMO372vS/Ya7Bl/uT6F6oEOylRpS+GmLgKNdpzRvjDPs8xylMa2K7vn/ppgwaR7/aT
JdcnH5omuKLxRgGr7J7AfS0bpUrsV6eIl9ujdRMkBue0KMfEmOnyyrOq9zTasNsAov4exE4Xj+8X
rw0XtSAV1EsiqC65KWw5oLF6XlfYwkJNCPembl4flBf7tixxuKXnROQUWSYC7NFZFt16jFi12Jpx
Ivpy+QWg5MjrLRE8kJb2iT7D7yG8MjlgZjmMJoBulhfmWGJPGuEN7ThvZr6gmXShhAeBHEauwV23
SU1S6hOdHMUn4ijk7GMbZDoOWsT3DNoVJ0mcGfeFjpYQRIFvizE6PyPds+VO0NFG1gYBKrPkuUzA
4PRU2MkLP7wwjukI89oOSZVvTanOvSU3jNymt9uK6K2KKHEyExdIzfXNkaJs6l7xml7a+0/JLrCe
ps6FxtstgDEiMiTFv4ySnMYaLi+VBscyjhj0EJ4Ud5UPnatBFY8PWiwY7SRVZpTMDLjcEgD8Cmwg
t0OXLuAbRVLk3hat/ncqyiVG6X/wfwcTcU3YzWR7hE42MZdWpg31QF0LSvmmVa8vA5E9rWOcHOIc
Dw1Ywr60aGL+KLAB5IGsuSOlVlGn0xh2gZzaa90fYtMIxxiuYcYX/qWH9n8Sz3aFycJAa3+JtqHc
jQ1LSGQz/T5vdNj3JW47MObFUv+SRA7bgoX+vV7EF7RGMTqTJCbF2kMzJik/7FLumkb2aen2A/z6
PdzSy4fQzv3xeqEu4tYRLcEXDrq4QfelX4Ee/IqSw2zxKcZgnd6l8AblZAjVH9FYL7pGh1cNnT9n
38T1s2VnYMtqxDfHZ5ZTlwvi3cWU22G/HF9XetQOI6SM7cZr6PdUUukIk98vTOhR2hu43DTbtAJS
CqG1hG62rh9JCYRfJQNF8IXJHOtgdVijhWoCqLAOhfGvigBQVULHZzUBygz8/5ArBVdwRxWpXw4j
4qsDItoxXS3vO5VSAOC8j/k41Ff6p346qUPj/SPtOrQa0uvEG4ZawvQCzJnqlS/wlHeFSUybFmVi
LNdQ4L8Z6qOg8YUv6BNa50iqqPgw6yqafoo7yDDIyIZn1A3z8qhYG5RibP3FdEakqORGyZIiRNQb
cu+suxadMfI6YiFcHFATyRN51NRiloPM/e3I9weL7vQe9Lu8v29WxsDI2Yv5m/1ZQCbjZdgB6SKO
KRY9VitsYzm8dEWK+MGLTpFXqGY0SfbALpVb0PykwFHpwJpZqdgt2g1Cakc0OISr7KRILVhRTVB5
OkdVHAOtzmF5wS5OP5QKZso9YUssEUIGBUAxT+Nk2Q81QTkdAhZGmfpJ/axXE17Yhs5Qz9GhvMRa
OZuxmD3F6EFrmbXAK2FLnHWlBeS7NhZ659QW38MEHCevbI9gyn454dTveviI456SvU6aJ1dsDFjI
REA8lr4jET+0n5UfFuDa5h16h/dUJ3QAZxbofvhoT8vOBMswgsyfJ1b85xk8X90qlxKfUrWU4dfy
boHH/3b0Y8rs7QXyNd1wdE/5gOUoiBNwNpFIXSc9NBhk12VFT38jPK2o5pqPT1DsTM97rCez0/Zm
KOeJDNEiyD0IXrecoebZdzFEesZU5xgsGCWE8zgVGaCdRVYbNa8YqXrLu7orfY5CbfrQlZMtANTv
FAdUzKGUK3RqIR4OS0YHbMP5AhYVlUDWrfxaAuhJHFVfq9KGjsd7yXVADoHcmPwcSK/f+m5c+m7L
BNBkZ+CdiGSeJME/4nBz8fYqwHv72Odlz3eLW12l1GSg8J8L7/Ew+rM/OeupeTb3YCJDUaTi1CPP
OwC1pdYw/vOZkgfdNm2OpNUeU1U7cEIIJU6MhfkdjUa+DaysPzm8+te84heymcejLiybswXMRLOV
VPe8MvH/GRsxVsqjF1BSrdGZAE/MRHcjj9MDpix3cpEnrGg1POi1aYNai28sOvKMMYmxxRJiS8Oj
uqvBO+dFymdSWD4PMmP+DPuMvyaPSelT4OqL3hnFzCB06a0A5BE4aANtvfB3kkp+M2gygeOveW73
gPMXPN6Dc69rtUPKtpZfrVJAd2rKSR7hLNVoyQGHaKF5mrZti8UhMT1Ql9SpyzN2q+IltaQKUdpr
ou68eP7/CiayLGgzJpzEcZT0yw6lTVimVzWxAipwUVYUqg2o/cIeQbM48/s1pU0ndBb3yRqP217g
6sNM2n2xGKgNf/gX90yh+tyvT3lffa/yeeXgPgIyphOC97mhgAkCovenKohqS/BLRBZoaP8QqKw3
yJHEmWVlY+4XI1oprSl8xkVwrp0ZfsmoYtVt8Nkl6W03dlNZosOwV5DF3FYx4QCMAJzrvpLvo5dM
8T5JDhsNtgYco6wWIpZlElBVqrPfW++/8Nlq9wyG70FeZDF4BsXn3RYCJGtptmnWx4uTvCSub5ua
A6EEgRvG0WCctgAyEEr4wp9/n4GtKKZCZYGSDzNipn/oGLilfoNrjQGM56lPEhp/9BwniuYeejNw
aPmJr6hK4miM+zlfrovTc5aA4MC6Bz9nKLwbuY11uvmMD6nJYUm0phSff8+3yh3WUWwzcGXoVEEd
bhynDUyA27QHSY0AnjUzrfTHuuSW8ThA5exiWoOKEaaVwL8Fx0u0okKE4BE6szaTvSn99onlOeg2
cWZ/wN6ty4etzl029BEtmH2gWRDdLQHgA4DmgRPB/Om12YMTKf32LC6xujcD3IU09s0mJDjRZ8zK
ePtXPIX133Tv2rjmki4DUIDt7wZXJDrDLR7Jn3bGVfoi4tnFP8ctoxCk2o1snTCR7daJ/f/L1C//
CEwplwJAHlCaGZryXngEFfDZ5t5EVyJWWBN+FLgZjvYHHqXhXLSde/OPTFe/2eQLEbKg0k5jaQXh
NUzP7ofPj/DRGHOpa55Z70+obF4H2lOk+aLQrEkM97kO2S+9/8fWL9p+P/2j+uHqPkoZhVHfJ0qi
ri8YrzsAj69MNXXxwWp784m0UIo5FRUWj1b1WCiM1urcEGCfPD8kRGqZF4VyguDbXLt6W1G2Kq4W
C9ijqX4SomYZy0JZhpTo5SurXEKYfBbQ7/jlnuDbRcfDVil6x6qVuxyE2ihEKguu8iDK9slQGUjQ
oG3/9bPpB7PFpu4tnY8egPVNYvYRDnMZwtFfsGO4QXtZ0ioBueqL9jTJMi/C+5Jh2g38nKCHAlPe
4nTFqeWFY43blZ3Qop21NSSh6uHZGU9eFlAsBKYCfzSi0LpWtSD/tPPD4czlNJ3sVtO/4ahZdUiz
kuT5kq4xX9MPpodKLoSKs96OlpczU8bLJaE8DfREmf3esZ0Kl1ohfRrCPxSyb+uILOZYs7GIMTcs
7cfppU8L7S+GEzM8o176MYMIB3GjNb6n2jFVW0xn96vvJvs4TmNBfuE2qjng7E+KOkYZcO0IfPpK
XmOOzlr7SXUnra9mtPdIcNax1wGXmcmmUzBKgHxYPgfyHgYgKXbrcAL5KlWGTL9uqe2IyExAOLUV
uWdOsm7Ua6Q4Kp7HQGXy4B+Pqe/bWL+sNau4eJlN8OYCL15ptE4bsWM/ao1lT3ra+c+++CGTZybC
GMOralp38IQGR3CR+ni6uHCe9aLvQkT5NMhQXgqgSOGGVakrl3njXZrZfVrqjr+9AlJlw1FjSM6o
B7o724Rx1OHeWSz4qEfVxoUb8TB7tBULT+C7EL2tAzNt61+ED6FSY3uJXO5nu52PoZSqawu7Ge9o
4jPzjRIGMJ91Ak9Tx7+xyM65FIzwSfBxLii3hGzVslRqEA24XnxhkPC9DXVtrA++bQUiK1nrpcnO
lSoCfbo9R6rvvw0adG53Iix7073PMjSIPCm6h1ZhWEmynNM+n7iY1WPR4oCyy4Hgu2bNu0pEC5ne
afmbX2aul7/5DYoHvohZ+gX+tPPG2OFXYnW2uDuZ148XQh/B2ZREqF6OkNKNFxJzoF4P+yUII9Ar
iJWacrpqwyPtRL4tuEahNIu3lnxQqym3rd6mnVlTPU5A0NKgo48q4h6CIB00arB6/lUJhgbYEvkr
IbCJDvbj8xF3oIkDo6NsZ//yn6+LwBYWcGcvPMJbv2gkepaHvjYDo64OSiCjqQfKP6DKLoWLsqPd
gwl8mTIN62GNeYNekwoH4PNiKRF3TcMobVIjHYEKQsRp4hjbL3wjFONwxxhYmGqAagoSybP5Yo5g
B4PFX6n5/3Dk2lLCQoYRn5+mVTdbSNmrAgaXiOHSR2zHcP7iyoR8zRhXd+hStPdiohvRQK3V4qk4
PLka0ped7DeqNB20X6Pj7qfpw6FI1u7jZXEbMc2GBt0xBalH/mU4bxbgmvxK8t2vZjkVepiB60oj
GLi+ReTpPVlDMuGteETwq3aQv7TNna0U2eIxqFp4ujj0CcPEd1pwqUIYOxL4/7bzYNXTDm0rA9Bc
/3AFyl/aiBSjfNzAOKsiaq3rrJ9a/yKaV1IL/SsBnEucGJZb4qtzKvlO916rHCrRx+vy+sShZO2y
iqiT4atdVKicIWcC7GvjgMPqWkkCJ9dKi4Fql1AoEyOVWNGIxLZA3nrfqGT4ojP0016XVAq5nNN0
kERFjk11SBIeK3jrSOIn/4Ks31DiX8I9ObsmdsSxIf9j8Ndfo0HK1D2jVhrKBVkz5hQz1HtDNlNQ
p+9Q+tB3P5evjKXxF/miJWxnyRtVU3BqzOJWe35kgHXryx5JbdWH6YZFgSmxvBsM9Sf45Zwzt7aT
N7Kdum3uMrZ6Jrq+sm8t/4UKvN8ZJ+8cfFeQnrNT2kphrCQvu+Xh7dcgXPjZsiU0myMdzPZDXTHh
dpaKAgEeO0bLZWwLsnq4Nq41SEVPI71Hk58j1nrmwqW/QEd5+FmlPXjMIXtf0YCX5rxdsH4YY6OG
f7oiu5ViUrK1aO5oouYszlI5rV55OUcGLZb/cq+peM4D3wXeZYOhLzFefkfOUhw2nvPkKqosZiWa
MWDTmU4xZOrBxUgH6v++PUW+iVkgDFi6wii1rNtPn9mbadiUfwEg1s1UuTu+WeCIyJsyLJ2ddh2D
eH62TkduFQomh3XbpGQlXwXBSZv32i836DOWzvZ5uNFjodAu8B4Q4iRRi4IwTQzzn584NYnHuy1N
nnV/2igZfBFlly5EARFnNGfc25vO2dvcogdCFn0iW4W11bec2RD32PH+MLVbFgYRwf7b7AD+0Lgq
gROqIIjYIyz1V90LOWXGMgi77BYMa/pltQRVssqxLCR3YrHnt0ngesanQCAR+twnPrOOIFXg2u7K
+c/e9zWQmr7hv1CVOPvNh3rJOBU4op4Y1ZrqA5UHOKTFWWkhmGgFqANDiUacIpErPTuHnhxNmTWM
g8VO4OrTktz98lWZGOF5xIh/ELwbHP/BBLcaHTq3lH2nXmdBURaiM0nEtJyPlMqupsOIhiJuWRAX
92DY4J/uECKHugkBzpG01Xsda8NuY0AUVbPgAcfOpqf9dsOZ10Sm4c6Aztw8s/Zad5imK13dR0Wd
6JBvnPiqyhttYJ71qRXJrqjmw+NzaDShtP4QZJbvMbhiFfubo6XHRzgBHpOcPcWoTx4422PNXP+o
R+KUokhuLoTMgMksjjQcFiBOigEe3kdEE4JPcjxBJT8o1nq05VM0bLd0FiFavQPKORkIZ4nJV7g5
+4TtLFOPyEV9mYGNzJtnkdU1bz8pCevlGLvuXZ8fDr0IA/pkBi4OVEHhd09FaGrW01jVgtfc30YB
AEkfiu6dTl+5kYe48OTpYdJvjZQLwjkEFHr91tyBfKUjth4dH6HrZAb6RVatgeJ0I9N9tE0mpnpy
3i3MWm3M/6oq23RW2w9FtWes+WUmNGW2B/g84WF9GDtUcmQ3Awa6rXXEvEQphQWC0PHSZt8zHheG
3EthQEODeF+4Lp+IBoKXgDqqxi7S67c91HxlNR4Nax1xF8m0BJyrMrdfBVW1t12gcuyLqHTRWj42
0pZF+nG+V+HvcQ+DEaaRMswHRGOIcYPHvGcaHV2JhmzzzzwfMHK+eLCw4enm7hfTEbuz1Kf49BQQ
x3//vkTMU288qiu5tsRoV63xPSeUWWwKhgBL30u8t+FFYfqah3zwhS0pbpBWa4qXhzSmrW7yTey5
5C2rB0jpD/c9uUZsP2CeouPhNew8AT1m9MI53ixv4+wvxzdxqsAleXwwdJFd2c5c6sJgZ9ytYCDd
Vp3FjgffDe3cU9z1cCnWfqHT/xeJJ9dOKi/y+HW0uln752Krzzuum39BuWD4p5ihw1BnzMs5NbS4
Ct2goYNy1aEqPqrzznOkvu41eg779GDYTJhK2M8CezuDJ2zsVbA/ne5caclnhkjigOVXj1nvpwvW
z4NNRQRNqCcLA0pj7wJ35GMJcuYk/NdOw9YjV4sSsBMzdcohEhqRc87+rpuM6O1mCHHP9/DDS1ki
UWSt9+AopWEGhuB29pJWdLjM1SoVale19t8ea9py6TJ6Qcz/hocXSOsir7PxY+7AwhOiCybLciau
r5blW3fSfNoW8u0gZqSP/nY+s8DVrQ0No/a1jAKqp0+7vtpcwBXIrumC8k50vXIVAmkzCeDZRnEs
RpdzHnLCw4lr360KTutNwlC99BF2my0f2jciwLO/364fjxldVUFEh/HH+zmIonNAB0rkYAKLgAJY
yDLBWnBaehiNFNzXAjGd4HDTJQZAHQaa/q6mgFE7wOHknA8EMaJQVwB8F12U09ZxEvT9B1Rr6RUU
XAICaST2xlxNcov4f+jEYNB5HNMufwrnvWdenWkFiYHNsqbsW9rO0ihE3ZxU9IO+sygDWVaAOT9X
XBjATtA3gcJxWwkt4nMO/oDpe2BWWx8CqUAUlBiRDVUQTJUlFXPVBeC15iaErsWEZOUEnrCSXrsL
x6gC+fZ7SHZFOUCMfReQ1Va6NUAkZ/00yjrrlLxHfi7MBKot+DYuKmcDSNxpgWoql/cMZpLkR9EE
mNes2zKM1B0guE6kdyY8uvASK2zgBLcfsE8EhsVYI5Pwf+0Yu1C0kjLkaC/wi4HwUsQ/3wL99lmy
R/RuDf7v2hSPES1oJWmHrdxkuX8giK7xCXcI6QpnbxXF/nt/bU9AX3gWobL2qgZzcFO3j0dw+Mjf
QUYr7v0kyl8D/Ma+i1bTepWtOrize5HPZqK5DUTA7+EOSOeels8pGndKEyrWIylWvYjpzlU3N0mo
IwZIYvp4Og1s0YwtaE8Wr87Ydl1rwRKUiudl3LcIkCaCQyzDrfYYtVW2lfR8XRxoq1MvmhKF0y4+
c91mvU13U6VpBe38YbsEm8gQO5MGqLAGi81N72o4I4U0q3I5Kb5Zr5ew4QfMTNMyHX+L3iSVkRqu
AfcaFQ+cLkPqBiNzhRB7XnCO6x4/y/2GjUOB8davKmKqye+yyUeGEj+/xN12uOlh4xsR76qMy8VZ
YdtV3UHjQmI0F4N1kr3gueFEPFgf23OJOtIqPnYBc72H8qk0fjltgRxK/YAj3n9hatqcoxXXAbjO
8XOtNfzeon21AGeT9jPmCktmR32EC+pxyhobJoTev44UTHe8Xj4lCoDBk+qXd4firM9AlW/HTSku
owAxIZkyJjvY0AKkg83xiRwF6Ul0ErD8DoaMuH+abzTz3RvRSplIrpwbbH5PHrU6PKD1WLvqfwuG
sWrX94r4Y2czy2P4Y10twn3fANsXkPAzZ61TdOXQXAEUOFugveXs/v6KpCdhdmVgQdSd5H9FF2XC
b6XkU2J/7sxiyuhty4K/xwyY0UquZT59lYShk24aOeT+qJdCMGSSMUrHzPVydKGLHTFq05BgZHtA
g+lootc0bdPzcKopHn919xK8J2vdiovL2UGzbxmABDC5NHFdJSZlOOoCzC7YA3RdhK9tREcgw4Ec
xpab/eKh/wA3od2o+KwgQgTGf2G7TAxidv8sOms6J/Ci1aLiXKbRY02peCP0wDprEX5jXa6oUMas
ZvoqoLERZF9LzyUH4dqLQyhgms5zON7ixv0gqIb2yqgE99W+zHXWlH32O/vofouDvbsAoNMpUNO5
JxYh9fTTsYXG/C/qTnlrTt6JkHeJ601DN1QgiN3drY5xt807hSb1dz4s0qswkw2r0++axdyKOnyl
okQRm/N1ykjcgZpqsr03RoBnnf2delwrNKsLO+J0vgqPNSpiC9a+mqxHfS8vX65CJw7z5Y/EJKCO
7FKl7qB3c53JoNQjO/8HfdRRW3aGC2xURNer+stf5UMYdYu+6X1DQDgR0FmoPXWFd6UH6yKlPHfB
sxrc9kxcOhvMWoo83Iy2jICQ+OlSFcdFejlJbTaZGOIO1UI7sJYowEDUXVNEbKfTNFfELLu2DVJH
mTEAaERRCfo9FoNBHzdpVe54kQoV4cNZrhZRUWeBjo5J7cgX9jqZt3gQPqC529gJoX0ovxh9pQNJ
Dt+3qPy+FC1r/trmzkWK/Uw1F7j+VJ+G0Lu6BS4lQ/Ol3E/JuwbMqkCRC2WttLZ00rJ+iv2//bg0
Wb4zi65/K4Wlma02T4LWjg5GxAY0nqBMxC+ESGVbJw4r3uYep1WsD4/6qo4U5m0jw3DsFNqliru1
+1Sl0HBxZizcBS4OsStGIdI5bdKcg7MWjqoPN+GY587YRVsDuYRutsKHrEoyMRCYpTABNHRNQ3jm
CXoZnM8iphcVe0vZpSjqoEqziIgJc95lZQVFyIkP3yGfcjYrIJJr/FvfzhQlWcxEEMnBVEMK7op7
+MCthbsZSq2Z1uUKBklQX02rn4BFwdvvzjXQ35vYEs5BmUK41P5UHATKVlDrTIP6YXvCfYdW63EL
vM97+Y4Tao5/FbnNfaGeeV20O1vFgz/rDumGIhrOU+HkfbCJNO7Nc1JuS6XcTc1DEOlvbJY57W38
bFlPDvYq0cRgUdx5Ti2jVAO2oSFbV+4cp7dMVOruulfR/3Dwbfx2vGjlTS+syZybcuIrWuVMr2nP
E6kkzTraJR5onLbvy+shQwDeU4qIlhB4uTRIH6in1GOnMGCMdNJnTdxQxiGMong6b9OQlFbytD1a
QXlBDEWDww71hFMXXW6q3rSeR2NP5QqqL+eAkyR232zxtJyCcOZ/3n5nFdMnpdX7DF3ckQ1TqSUn
59/foz9XA23iDo7oiK7lERCrEf9NeBwAgiwFauv6Qhwf4lJ5v8Hnal4R25x1eJ0lFUFPrsBBXAyV
SzRbE9YpiP8irZ0cquSMoH04eK8rqO5EaKYZIXMPw1uoEGLTHVy0W+4OE3VEYTov/XwjWMn7XKPe
bEYB+a8fGSbsADGRMlqsd2JTTBX5IDTvSlz6INnOaoROkPx5mIUmE+6/yqu+aRxRbjNY+h9EfOBk
8qVk1EEDQDt3XWt4unD5CzWrShtPp0jWgF7M+JedJVpsDeTIHDnuzC5ALKRBGRDP1S8fc1hHDGCR
Nj76sct+QlkvUx9gbKzw9xB+El09xczUswmn36BlHG/8I3LsOs4su9LcOoF464s96ZYL0Is5csqP
J2ja+iB1kTku2kuquGr9kgdwudrzRynnIc6fjRbCn8O/9QK75UvU2s0JWyNGFwuwF5Wblp4EFv+U
/FG1zDHkPQMQ7JDE7ZLKtxMRkhvXOoqqVw/79XK9lKRUDmXih//juP359Pdiiju0tCoyF+y1leal
wmKKC87rgqXArZSWo3PI91aUCO6Tgv/L6ApdeM5WjjUABx+hJS+mrkUrMN7YpR+APcLNALXtQr56
6Y7UTFjpPABm6rbRIVB23an3pG5B9F73vu3glpgpMD1kKOZvv61YMFfeNURrxHW9A87FKnwZV7kv
LNi5DVeCNRFl4vyA0HH9ovqxxpKd55cYM6rwiIEni7UwUjaEXCUS6qF32KTtMg2dPtt4jlVH/2fd
iT+FS/9qv1m7pxD0tfM6p2pNWtfkAOydVBwBpue+VufETktJM7lZ4XYw7QfX6Tcqs3MyHN7KyHIT
c6zfQvB3yROf7+FzcsWeLZ5yB3FG0Ghyx62SWccds9Vyx3wkGxzSm1EXQ+PBuE13hjJg9IXRCM/x
5bcVoG6thU2KqX6M5zAmP3hGCn42jpEtfajpT1T60rqYKyJj8b/R91xpc38P2v9PRyiqWCQPqJWA
LDTZfdWMyIYeS54/hDI7zy0TCebIRqvbetVdAZCNEbmJHXMq52XYBe9KhqN8mPUkC/47gG0ZsLwh
VVo6qLElA4JgJZgP1h4ZnPwGCNwOdmPxWM3RzrnlpPuC0pmNBr39RfyFElXVRVYQRADY2cQs4a0E
Qgx3UCwCIaSiKSlmktsEcfVOrQSKaw4SDjkYGftQJILGlAoxBo0EAbCeeU52A0qbHOYO0hEU8B7v
/j47UnibXtmnRLdWbGw3KIJHBJ3P47+QrIc42egcfaPrc/6/1YpZY8xcPqCxhL9VBc4R6rftFZg6
N/OQCgiAxnsgRIrYUpw+40bjHmimAYcBwdrFKhE/oOVeUtuG4aQQfFDTSi2ZXezBpWJq/E0qgErv
lMe8AWuTVQCMt7dv4kZuW8YkS5BK2GrBY0BLOIagv1K4IEjaiT5amFX3WhvwcEreFWTr8E0rX7Dh
Y53X6JkdVN/LYsLeO63OhsaYQ8HkQ4YQEFXx94H8CnDO8wD+ddQ2w+yN5R0GDZOCV6iMaWtQBzkO
jg4/+RYB8zt5x9uafSVcCWI2mQJ+yfKiymYG9ZoU9cUk4dJACvodnZrRN3FS6T3V7OVTAsX/Uwng
c17Tz82bK78pp3GtyC5UY/dhkUjTkUc+0x/yB7Zrd+RsXqgAec3ZtYlJ1LTEQTYZDedPg8xOTNE6
WdX/RSdJreyRSl6mslOvIU4mfamJwLmltvaK7WhEIe9kCNqvrS3FdSkqem0PUnV6Vam1A4r5IL/x
SSBzm0M4WK8P9YvOejrL4AxAkxTN6zrQsl9jj0zeVXTzukrX73+cLfP5tRRT6H+nIyWyEeCP1VaF
NGFL5ta7dtv2SyeBOKWosXWhTbS9aYpQlfOC5w1rieklvk+VzboXy66YRP8AS6qAAcjIUx2hErN8
kGOt7Ct2NouDf2pekDW/PeGPKetxhdnxtsFK4jE0ZpUFXmSPUZm7rkcg8OGwZcZZulCvuapheY1n
AWmeT0NmCIsZxzmbEESkkluja0XsGeFTNueEjI14GvYkyNKkAb/+svk7/U7qkbNpmSM+rAyBsam5
zHdLqyVUR2vxuKhx+ex/l9M7egyXikvM8dF0KR4C4pgF4vxUsvI2/dzzVXZRfyppq3Rlqj8nEi8S
MhPFOYmEhOZTple/qIBxVq01KcC6PN7D4yy3KAaWTdC+c6693vKv98iGGUo3QiBQSOvlP1ePIbNS
+zaenMa/yTEhSGqEjPkIP6dmlfxt93KPSAP5pnbf+bc3RTK8WRx9o8S1cRKpcU4E1PqoGpmIRXql
wqSrfFIjFDBXTiEow5Te5B/WquUolb7cefA87ol71bA72FEmGEL37yuB3RQMqfNPhcgcWr/GhHsU
1PTwP2HdXNdI/mh9X30XzdLyCUbMpcgAVJ/Pz5BD3oJAnmTURo2FhwXGzz4xiUolkXiicRWB4xlN
Q53d/J5SPHahscYuGDFcshgURXXXP1aIcul7ZjjOjpYGlf39DiiQ7eDJUC92vqGagVYH/tkDDwl4
8d5LV75JwRk2ni0aAMJegb/5ymGcehWOozFkhmaR54IAMjAJifujnHaIsVskMA6wXj1YxvTy270B
7rSxiLalKPDBurXXB4He8ri6M/ev87odzw5QzGup3NzjbgrIMa8Q8LZJGrLKnzdpoytMlXZfJSJH
sDMdzVhMt2azQ4U+TKOi2TSYByQ4f06CZxTJynQp+Xuv3Prx9wQo+Sh6MVoHCLJkJW2uLUMgKUf6
Ofu4MJmO43SwrXoStOSDYza+mxe2BzjzrdxE+1N4Uxt2T4yOQnsNgkDF87BOUR1EsSMDi+CO1XxI
B3Q/n9nE/zZjUB6JZAh6V2q7nwNGQvzPOHyNsiAmkqaq/P2Akur0Jk9LF5ASpNUmTsIPoDxTF6TV
n6yf1GTDHAsaIE6PUxnuaxTQPyCA08jTJNd5/cz0H7iE9ZKznRoCMXyQ1nI+6Wt5GRbB7Wj/6cD8
MFopEzyzWp4aKFRLJbV3PDsSYm47hAOv5slUTvupeGfDsQyZ/95h8VztMFNzCvn+4jQRWHndeqYo
e1lckVo4EbVVaRy49Ao7qHs6KFdAFxnwA/koj1LAoq8wzY6k9VpQD9NraX1Q5NhrGFL9urGFE0Lh
q5bQ29uFXQ2eDCS0b2+oiZorycFMPkxkvNyfDy6DimEh/aIbBskm0UPy+E8t4jZA7UfscJYYpK+8
ZXfqKtCQXqbPqifpOaKk8lNB1C0Ry59zYr/bf30hRdjvlzvds/+1siciKCEb/Rxo4oSRg9S7zglB
4zE7AiSGJ4M5yhC353/xijnP7pB+/LZ5+ywvhW31fIVpBMpKVEXv13l469m+sXU12tuZJ3BTeRtP
4DWbSaT8Y6xb3rv5+gwlcbYMvGaJKI00QpuVurcrIUZeeiph8MeVjn8U9evW2/O/N7V7EuTu457X
NH6NWVm3DvzRDvn9zoPqlGV8bPiiJKJjGZ1rywoiXMRaBGxDlUJMhwcIfXqcALJw07PVElDHpQ9+
UPfOPjjBV75LaQvOcAVIZEHg4+w4TxtDCiHqSBMNjYclEvihaO6fV/07gryrCazUO3JLziPu2hkc
rVWrfd+dkHukMfnAmcedqPH5l0hylX9c/cpP2A8/UOfegYGK4niVuJ62eq6hetdyN8pP3vCiK0dV
+a2jZWlSZzTZSV03tFF6QepA+tUp3FrtXj1FVPstdGZyVBd4zv0denbnPGA0orZDvH3mn3kHbP9a
AhTfWtEOCREwikYAhiGvL3Hh+GGVG8xRi58QXFpHFWUNq/KHI8uviPsKUSyYz3zF0GakHLCPvtMp
JtjQk/MWd/kwAaUJalhvDD+RzfbKyfFlsz12gJI5QqY91HOR6G8YxxCQZT31Nj8p/GlKIhYYq7qE
+79EOp6+2gfjrGQ4L5DwG2N7XORcufOzOpPoCS6G93YDc8dh9f+SM5rDZOJvLcNYeIku+QoDBq2G
KDL2XVfWFy8hY9GwN3KMMjBBNoEFMSh0MjLKI+6y3oayGPn/rAI1j+np+AWse068Aos0mVYrqhIW
jhCuyUCxAiM/TFf30J44GqDsImVYygHzytyhgPwHF6jom9/mR45EwB28z9U3FWHLhMLQUR4kCLsH
OEUWfTcMds/zW1U1GY2IFxdVDHyCB06A2dm4yoDawgrXrobWyYe02k7gu0mZgq7ncbi2k5ANmRxY
CjcssLZiwJdvET+BU+GeRIGChyz+VJk6eVUtf17dUyToJk9ZoCac22UMwJlDzQShJ9nLiRaq+bZl
q9q5WxqcvCOHaYPOjhlXXJ40JT1/xb+wubA2sZ+xfBB1x/8XWCHe8JfKznx9Y/tpPj4l+8pW9ZL9
X8asDg/rRjkug9k5JQ4jFYdiQXJez7f/8TMfqTCGZyz+p8GbvuUIVQAt/mr1qYWNm0sKkDkw1snB
8Bb7KY22WM12aPMAAKXWUOxwK8WmqKtI6dtbnXzVp+wIImeiWGHhT8H78b065uMBkqvOH1zIM1KR
Syi2f4TI3aGqjVwLiF1pIeBNagMjH5Lz+FaefzV9tJjD9qsz+J57KoOUpvk4AbrML0WITa6Stj3Z
PClBkPieSUT7byfo2dbWUWh4OI+NbUwChWNpvHrmVXeKdwDIiqx9KkIE+wL8gJY5RaHuJISgNgr2
enmOfN4wqhBQCWCc0AFVJZf0lnxvPSyE2U0LYuPOsDRLD2WeJRhQH6RHPCASgghl5kUqfqTGIZVT
zl/ls1fO9kUSysih1FrPp+Ty2GTV9w/6TnRuGiV5HluQiYjHrZAO9st/NxELgX/JNRztl83zVZMM
dBGTM2jmPXIo+U0XOR90TLs7GFuZ6Dyv9Aj/iJkO25o7yk4rSxO39dwswYG623J4iMbT08cVpLrn
G92cIB8Z4mv0H2siNpQ3BTSa/yQ0ZMsFdrlV3mNWOJ4DhVjk48WpxP3nzXK2ZYpKsn4hxnMWPo9q
CZdpEjeYcjK/qy/FkgMv+Er9aLPY7/ZBAztVu3qB+px0LpgYv27AvN97UR5VXVlMdD/NyxIdZcIx
sjXhgS3J6Gh9OzG1Pa4SwSmG0KHwIulL2snnJZMwiDkQLDEHXy14ypTinE4zYho5+oR7p4NQ+Awn
T8sB23B8FtF7f1udNvTxbE30V+2Su9a+Pzpns1FcCx6OeWQLRGvlf9K6DNjWP1iu1PHdfoGF5nB1
yuzficbU603hlYp0bA95voJnRF25RwIGh4AH3c1JCQHbD7Epd74IxolApe6CGUGVmuhOgsmNShL+
V91772rhmkwy9c91MjJ+Nj0/MeUnrIHQrPhczblrRE/8vyZvmN6MKanpPPA+2s0RqJmziLPChww2
HBD8nwQ8whTP4mzfMNGV3U4eeMS9F0TVk6jJl4+oWJ6OW5JpuZxUww1yUMxAbbxdmtfriJmq3h0m
oINkUsPhR3GLPha1HccD019VijZnphejHk9ZKE4kogvko4b9GrxnWRJxhFoJ/+7GWw+IKpFo0P/c
5laY0jjYTwWP8oDL+bWHLbnuLGfnnldlYiUU8esU0qHiHVwNQNdY6SDEefcKDhDDSF6IM+A6EtAQ
0xmVAbkJcOxobb5RaowBmrwRli7vNGlluwfdYyX8MKRXCoRSlmDqYLMI8WaWDjj5Y7gKQgG6Zecj
z+qRDkv4FFNXd5+RP2PBEpVx7/C9NY77FKEHCSR2HpTF2EfhYQPAU7L/Cy2yAekvPkyEY5YH9J0K
kJgym94Z7y7X71kHwgBwlZzuzPArOpX5i4akquBdCW03OK1Bi3r5f+nkvWrrm3Kbh4olTqj1q/Iu
bN8z6Tt19oyMkiTOgCrk+CeL6m1pze9Zlo8BHUm8ItT3VhJo9Z/nHGY+QDIbNTHkKq5Q2FPJZixA
ob3qwklx67Lvx++0oOsoEgpgJj9RCI3FVfBwKF/HggoHEL6Et8vnjhHTjDlbg/FPLBhjqKSXOmjb
UtUY+/95xmz/jXO3TQBnK527HJSxe/s8b3J4OEvU4i4Yfeqt4ZlEoauLLu0qR+Ktw4q4PquzjmCw
owX4I9AKbgPtlMPFg8LBYDS/tbFX1R1ar+lMTNyIvoPGwkYD2Z0YZ5Q1/pkU0RRhfBZlkuM+8h17
mnmtKDsyK3Y2xL6jpbCcI2NliYPKBqRtjEo0cSMDuwkNezQ3rMSplHCPJojTPtUxRYj/BNTtCs8i
lVR3f5teN0daalFLAN2CGprSwLBvBPInbZAIPEm4S0WEl9bsVbk92zXVoeiepadmiJmlv3mbibRv
KgW/fGUNVo5gc1c4clJKx0jZwEoXM/i7CXgQePuQbtjv7Wxnzamhp+V4kEzPqBMdXxMQXsVzxS/Y
ndhlprDylnAtf2ABApPEgx2dJkrayXt4P3FpLVH1hRHS7FwXGKvKX4deWeB85W6ka3OuD6slN1FE
cqeuJvXt8udBGsU7EB1VNkoE2QLipyvgpKvjOJDfuisgl1IU5/blIQbz+QlDmuF10Ff8TJH42GQM
WdlZt7D5aTVsjooMbOoL9999RNvA7Vz6m5NPoMfLHeVna2kS5LBZZ3fj5vMWi76F73/TBZ2tWf2Y
1VNYz/ZX+FrOgH999JotbDGOAj4vxyuOPC1847JPodvxsD1NyXE29mDx8dy4Lbf9V1jiVTIIRVm5
l7iVQN9eiPh/wmACnUuhGlMpaCmGO9CfHYcyes9AoGbw+dyHCfH9zpFX4UiBcahfdMG6cLdh77qD
vIPumxf9XYG7RUhMsLvsPWmDi0hZ2OX5M4tszwwJ2CBkmdXDdpRky0gK5xVhkkkcTIWa7p7vxdgg
/x+Oc5Lq9OeGye01kxNnm45HNR6CV0N4H0QokBzCUZxHyWtmtjkGV/43EQVVquBkbX/cUuPuDYLh
R7mwL8yCRw4W2+XFBj70nLbRCbkI7jsgweX6ltWmuudgClmz8cLNzcJXz2kTpFwwkRmnctr8Z8a3
Zd6BfgDd24bg+M6OoZP25EzYZt50T1xDdYl6RnnQ1luZ64SqrZ53cF0x2Y3HPL2dYnSphZtAfbq3
vVsrAHUXQhUyL1/1/oAs4WEQMMOou4bc4KjAL+AzpxNDgiyGoVlls3H32AKtNZrimyv2DQiwJvLK
QcwBo4+7tmwxDrin4U8sU+bYf2+5IIOu92o+ArgTXEPgwFfRBJ0VHQn+BcIb60gyZFzu26AWoMR+
VnFAA8mHXteMxMfPrrVa/R6bFHWKGKqVOjwiMK8C8gXH3n3xugL0BgOWim3YdNAO6h9CDJkzlSxF
yJxJjb/aXVXR6YcUdJbVEozjEzzSfcKy+rnLABcB1E9cPaGLS2BLIpBXx2XYIL3gOiIbFUsIuOSf
5g2ljmIbVMKpT6d04LSacBXDcwoCPIvFLRGPOHotoYscdpk0bkdMmDCbcK+mq0+a/MBMfbZftFHc
h9Y9x139NqALwgC1AttnE7ecJ2hw1hYALmlZpDlz3MHsnSBU9Txj74gJmyL9BelgwEDMB1PCrgQS
BHt7ABma14BFHZSDLgH9ZOPl+sOGHqra5JrWKqiYsHw6I93laz19XKgcxU2tRt0RcyV2HA8Xs+dO
5ECK0v6QUmkDvUKnPzgeiJZ6lhn9ugmL4dVwSorGHeLejicfPrTRWT7nj05k/jBUVWvBhuZdJfpm
h3VFNj/0WCOwMOKqPbYVo0dMfgmtYv9Qw4uV1CGK3xT5jrTRDL5b7JrrMmO6kV0ZyS23JI4XP6bX
NDoUkQb+KB2es2n0lUwluW4HJZWtFG7zyfvGcq85TmvKFiofmMbuZgDjEwdJ/bTp73jQ9W86DcW0
gV8L4v3YgIk4HhOUOpctYLWF1zBfWB2pE0fSMstEOef1Bx5/9RXncibafAkfS3Gx8OfhHZ+RxYU/
Yw/xk+z0mRp/xVA18RisRk2RA5ARfVDfIa9/2/xOFgn2QsTUSCO1vGuyHTBJbeT2bTF43aZPTb3P
TmsE9xj1g0AmRhAkQ03oR+B1kGgRxMydCUne/F0s3H9kIDT8wsbN7DA2dlsKb03F65SuIafsy2Gb
Uif0j+vsTq61UlBeAQxvPegkkvCFCIGW1mCBLrwyJFttt4sbly9ar9YjkdnP0viZBiqQ8o5tZzoB
8IVY3iMGUvq+4uZo0e7RGFXL48SC8vMJq3Jn0SkIcw3fSR6PzbtCQruXL2l8lKSOepEW8kwqFlu7
UJLltvlQ0mGuB/kef1n2fjR2gUuNnIFpVXo1LT5GSG8rr08lM6L41mlyAbevbpy6LUKgr5lnGw02
ydkJcSaja6NxERiFSg/LiEoTLhpGwLaSdF92BCCz9ntssi54PKvBXUKXhLJE551XH6OXrAkcu7JN
xRK3NTyW3amjN39OCtp0gZ7mCt7/9XTK9oh8mNMlT27SU4vBeVFsPLtiTrAYHwVvqeip+DvYsOQB
bS5Z5+2Vyj5xDLf3/PugVce+HGW3o5T+BAR48Zyfa9tmQpFrzYsApCHrIAv5cjTOlewb4zf07kta
o1AuAfoLD3UfRX0/0Lhk+8dmeNz9mZHIBFB0e0Po1SCV5E6ZUmljN5AZCUb4N0Ekauc/J0UZ/tcN
hsHaWlNRZ3niWoZk2hSEDlVFhqXLlZXYjZNmKyhzdt3sM3J+j+ZFjWZTANlYc7cVVx0Oo37IhNsu
1vmGSXgNvHGpfUeV/kylvxzxAhW1LXpVmXzQ6KmjEYpS4tOcaKfKa8XGIAJbPPZQPV7ReUntjSFG
qftpgeNo2XOs+ESskN12ChXD3Y0hNnWdtoPSrmunutCzrN2or3lJ6uCjRMXZYG0jc4eKx3T7OhNk
mXYUr1kqp0vK0/vTlfEiufqV56fk/kw3OE/PwZ26Ap1qDT5i21zz3rox3+IKrSqntmtUNc+QV+Ch
UhmbS0jxR/A4gHmwqtjAjo0TEX7ffWXqB+URdr4Sg5e6ktvaZ2bUdSx4hBkFtqub8GityQuQoj0k
D6ttdpVwAOevpwD8Nx3fTDl+ZzjsRxo6N+8MMzzcqJUcnpILOFYqTLbT7NnEzkk7j+4F0c/yICsu
oulUHj2VLAUrNwjQOtrNcs8U9iR/WfdMeDn2WlF0EPRUDmABHoQfZ/NHIsFnkMBJYGWdDupphz+j
79Jt7QEZIg41nXMQNwGKEapfLV4WQEx+toBNrMjyDCMyHD2jZrCQ/gZKIyMr707twMHgBGZo4//S
yy3bPL97O6ZbJ9SkM7wEO3Dy0D6wezV2EGfaqWibD2pOuqYv4EP9Z7PacOHsweV/u+r3ixBBzcnJ
jUnxUuSEMRdYZ2aTM+lMd8YITGwPd8xsxr9uqY1PWkvKCdMtdW028KXEYF3XdbNDNQXup++gOnkX
RTuAhUScHHUZB/x8Gq2nNihpkIBOdrWRkvPrvXwLcm189nZyYMUpBD5Iid+GMNwcSy2ZQxDJp62v
5aXeA6X/M/dFBJASTrVO+5ZD04BrFPTkT0KmoQiET3Bqxvkxxk9wbzgeoBUEXCUraBK+QvbnyVZv
rzVYQVqnYQka4tgvGedG9P/5vFHwNbO/2J3JSz2tdntbkmE47O1071NBY9WgC1/g9D0CJjNPN0/H
82Y/IkZn+KOwtelYqrOi9FgWMkHWZoK5MN1ifbpDPlTVB39SHjLVFzhsZgceEFA3T3ezSbjOdd6t
H+f+ZbXBJUXKqzdwA8OGbssqbXYiEHleV71GJA9aJnCHZXkUi+dmCqrvVPsgFQPrL5UV9RW+kr+P
kJ1V/zl/yZHkDpM/u65Rsiy9RxcDDMSwxNawa3ajuKpotW8WanTwP5Njsx25VTbMO7gvOA3+1fpl
fNW/bC0mq3P2Uk6GwQpBoxN3mGZq9q92iKoOuO2akhCjsvyygMmZM8NQexX1aI/Z1bha4H8pjvZx
89ovrQx2Qnr7t81hdRFc42rZ56g8Glp0lEQKneTcLuIAq6hheteayofrnkGWfkIklsifU5r8+cc2
wDwtH4tXIso+cHFba5wfA9v6XTsX/g6xhU7O+GHM89XINfcAdAJoILvJfBJDft/aHll1ECFhcoKn
dItCL69uwU2JTQhwTMipi7dEa43O1VxZuypqQn4rcolWoKQIxnk+L0gVzMUZAvaUZeNBeuMVsZdZ
Gwx/gSGaR4ez/LbWB+J7UuepP/cCgkm0WYogdjQ8r3xeK3hfg84iwGH+HThZ0gQVFJSR6G0oBum+
xKozL9KWKf/zvO7JtvxhZBLzXKnQfDGNIdb1W4Z3u9X2RHoGMCiM7GsyKXC7Q2povxfS8SLOWYJm
eUF1h+bZRNEJi81Iad8IdQp5vlfnEwxyPktb+sVRvnEifzuVnz3z7ZBDliq9HctxTE7A/jN3ID2V
PvNlDV0fKsmKzSQaCffPyMbkZu/OOTWsvwDtqAO4TQTJzHDPw41iz2+SrEfycRJTxyPX4rkAY6RC
4sFCWBtiJJrPBRwbke+9w4bFXbVRetW8GTbar7aSiTo7P8ItrybBAcOuHDBzzqTzwZ1t9mYpCSpl
LuaVeeUDWjaWbuoTh+gHFp3yZ0yhLLY5DP9FJQnppBoRwYuqcKFIzJZagxiFiDU5XYH098+q1hxV
kNRhKpw08Bc4lgkIuYAAcdCIpOYC1TyB+bJnIliV12hosc0Jtr+u82Xqk4prRyYHCYh9R+FjNkTt
AOy5mvNeWONul6AyqbhE5yRqYSltJjjDELm2qIqmu5hkiaxF/aD6yVBzk0usOIzqCNLsiW0xQ3pC
aJNnasEGDq7Bb5yAeiNvuFO5GgqtweaxchS9EPrgHHgp8dchfmLKAtFxkBA5KSPYudtaWzLMzKhs
28j3yDNl7hMMWPO9mWRtyRDOb2ZCAwDL2JOhnD9soMpFKvUDwe53f3tauu7pmS6MRgKjD7DJPs7T
MB2+XRcbnS9GBymoWo8wG/Mdusgq1drYiXWlxX+tNbkVJeduSTGnpcemwq8bpXdctRkFYO9xnGcO
9UFI3fCNIJFCS7F63nbG2ls5HQnHTSAv7jGK0KAxrI29dxCbZC6yIoA6Gs9Wf+pIExqu+RqtgfC1
iKPF3epwNrO11RS0soYhzh5O1cI0doJvzgfEGtsSwiqoNKsOAzLFwsDGOwty+b7AlPu3XxcGRA1B
BerUPqRaJh2GUGgIpPZUui7TbCzYUjd8j6EuaRA1KdwBrZXIIQizjCoXKEOJ1NDYrQI0yo4RPcRI
w4cCLoh9dXgBUv/L5Iqj22J5ambSqoice8mbuNkSJ21PsH/FKQe+uCkR0/VichOtuX9ltSVLITMC
IbJfOqjiPQcuL1utEUNXzEqT9TA7Q5NMP0OifboW7OuF28Bja5qlk8cUvLgPtS8rjSfQPX3wn/r4
WrAHgRIXGDHlb1bkWZHFNbnc7w8t9qCh6KrQacYPytiVeOwbA1W9CmQYUI8grnYNJQ5hQ1LMq6te
l+a6W47HlIPEpsyUHv/0zJ+ryToLtZ8P8edVvtLt5/iC2BBecLre5nURZpPdb7mBcqqpFIWPR6dK
EJb8zEtfGgy4CI2eQoHi1rFalRl46I3yl/fqp2D7FtBvwlJDOY0FjgNmqVkGE/3kz5rOx71Tzfxs
6yHKEX+7xQTa81pdPwGtwo6SGv8ZSkGalnITyni7TusVsj1rJLrS0ACMmd3I4YpjqWSgY8OhL0BK
4ykNVAYipiBFPQlfRoesy6+k1B/ktcUFU9P3k+8+ikymLlaminvAmdxeSGrtdsb4aKcBQB32TfPU
DdEsiaV0aiKB9wLZaRGxk39GXYBqhbviVC8+TxQIHkO8yxMHZfVjWp9D7g+FExb317FA3khOT6eh
kHIqJi5pESgvc4qbsU15f7Rpi2CrqTH3eQl6wcOZiubiYWiRSKpyk3ghP7PpZbaTRQv5ZbuKMV3e
nMSI1IWhesD9K/eBD1/aUm7lWKK06xWsL2rnYBr+i4sTQ+OZjiLPhGXsiOEcZsPIGojDbUA3Zk+Z
mpXs9z/SHmYRz48AO5/RUmVDllL51SJtY+5GFldm1lMEVE4TA2X6Aei2+HAPakngVdW8nNhBFqMg
KjAFTWOyXQaXiyOOjv0pJIEvT8NP+YhLK8vMrbx7IalZYVqlJZ6KCFSY8DE9ni9uVEZtvnDbm/DJ
f5mxfheX6JaHedynviwfGM5vMWXkHNU2pZmzWfW4Zn7vmfuv2bmpdLo4LqRYrrqTX8UZsjlPOlTI
5GDLa8pO+1gOUmYOxLsocKKX0pKTPxUKmMsI0EvwdkkTCb5SjWadvqVWKeZQlgSl6iJVEBGDp6qo
J/tjqc0IaANj7RjsQqgekJZPIuEuqfrvxTIY1kARy09c+C7Fb9kW31lXTJko2sKkQp7ZveyE0xSe
L+vvGNXfeH8BIXt+caFXnhOIdK/6MKXvoVFPUaVAV29BPSrsysvBZgnjLdcmwrm6uEx1k7N2LaRC
fmpryyMcMEw5eMn6O7oOmlVkkJQw0wn/4pHb9WNbap4IlnMpyh4umZA1GeauYhZPbU3AHahiinXL
ONUOiFKC+nkAmdG83L4gG8exfNcXagnX8uJvRif9bKw5H6P6AJNnAyROAlk3mfpSSGwyptBS50WZ
pxG+rR6kz1OqFWQ6aMuDq3Ks+8qFij4fenRo391nz0EJox7TLrAB9TjwuHMP/pDCxrvWrkWoH+Vq
i383pGVPI7TUAdEY3NKo88+xw21dBVaw6hB4hcn1i7nDz/KzkiI876kcVwePKjK4VDJ9NZpKeD/T
VMXzmv5BXCCkT/jM5/lIdcmorwkD61KDNh44mGj5f23yCThgwbsjz10CW6+N4qrzxBmWUImXCT+4
Vt8ZLz4YnGRw1fiZQX0OqFgTvmz0QThRzyC/PIUN96llUwBFuSq9/Tlq+HPcCW9U3wkiygruK6XE
cPUPJGglJObRyIHmgqg3/PG9oPXNgCPvKHiLUUsdMmrRJoYktyJ/TV9LyMQW34XRUiCZGI/30Wad
O2yrAlaSvanHGt4MPimFbh4dyYh4l5+ja3MYEZByuQNXjWkvl3P075r/CQ6/T4DBGqzL6LyU/hG4
B0LbGJatUU2gMsmdztyoWsGbYypu7rsmZdg+GtkLvKGLeWBU6JklecurePHE4fo2LsZn+AhWV3ca
5a99sN4QCx7TzXiWSF17nN8PXkjZi6DTfSOo7iYBcxIVE7srgvcw4VCP8VVf2Yshx7hGIs9xRCef
rZprGy3piCk4RQjNtuBHSK0l7kcMJSzc6uJmYrc5T/o+GOXdS1JM1NAm+mw3kmcaM6lur17rxq9w
n2hM4+H/rRncS+3Z/wFjjD8rvUdfQV5DPYzcgrtCgqfKeQCSzaM2lAmOl9QB5I9hxoYocPVwGqlw
kAvjBJGcGYG0y4ORoiSbJczV3WKwrIy5E2z9HbkB5TAxxeHP1aLkv5NaNdBjRyU4TiXaO4l0JHfZ
/oH+zhFYHea521f4PGSiwZJGltD9wWyrGP3Vp2DeUJiHDEFvlRpHvTVLZxNvCBoQl29De6KKiVBN
0Rz5xqMQkl4Nv1kSGLosSfrZOUO1KCn0wjI8cbUSglut1Zi6CwlVyDnGoUphTlktpNwhx3vITsx6
Q8r12HwNHrFM4Q8YhtDfrPChJTJw6biD+4GXwEOlJ4oEAgKAbOek/qf90FtYl1a+EOyEES9lp37N
sAA8WqPG79JVQBE0nqyQ5Jq0aSEp77FIjhrqHUFXDAiC0BX/9qEUt9vmqACi7cTWqWJP5qvxmPKu
ecsUQc6/b38QaqEJxrvz1MMatyAiPq71h/YsNZCtSJRY6YFhriHI9uJQ2vfclXgglb6FlJoCwEqF
TgWJdB5ltsDXwQJ+RyEW5iiybt2Hs52QMPDj7G42EEpBhcnep2ZqgyhpIXN8pbpgAIMQwT+A5pB4
50eIJMb4D8lIQjZwHmYtQ5Tx8beudP1oUXUjoPjgYcnj9CQ1cX6wwpsVouLFNOTk9VQRIjv1r/0j
BJwxymvWOb1q4df96dQYs2UsZpcM7ZLxBW/NFUT/U1m3MM9IKJ0q2UiL4RwsiDhUJBHXr9XEHpap
t36lFKJ1xSRb7Bb43sfhMkG6wBIMbEm8byopiipfJGbSUj7whwppQ6/DmxxmvDQd0qbUoi0ZD4OT
ogWUnIOdf3vaTxg8FwMjM3ti/QCZ4/NdX4WhvnnZDJ8Evwg16xasTr/cRjs5czFeXCvK0mDjk+tJ
53tWLDFVRyt1HivgsyaSs7TwfszkfbMGzxWVxknkmooYQfzw0JEtzmevsLQ2DYh0O4BRplKKMVMT
FuJh2fJLTiYtJv/D8AFev6eqLJEGdvR7rQzvPIBZyW1WufvVZVS9p5AoUBLSjW+PcYcOydLGy7Zo
Vjr7+YNCPwkHtv9dfQAS6P60xFcSJdX57DufrnjKu6lmo42jE58HT8ae4rCb/2BnS4+yGHYMfivS
yFzWLFRx6fpEm+dNDIXP1cDz01Iapsfg/e/ZIyClIfgmzMEg7gKRrPIOqo9p9Va8PHBz1BhCkv4+
N9QuIS3fzQezCB0Ie/UMPqbVqEqpYwvSPJR+RGo8nrsnR8kSQghg9rto1GhE+dKC2qozSl4szUGt
p9zW9VuImCqLChV4ddLfeNuiDXzHLc3CtXyBSBvYuZD9uP137Mr3qMnKl9q2ccSURP4Jche0ln2F
0HKbg58x625LblTWaWx5vLb0NfguA6jNdAU9lW9LZwVjywRnPL0n0J9/BN++yDK1XNuAMCqfOmSh
9g3Eomb14cpqFxsQigCzBPW9bCF/neGkaZSqhkWeQkSFgVZuJyKW5Lae0QqjmvhTE9rckZA6Awx4
GCZlULqP1hOFi8UgtrmNfqcJZehKa3/gvtkhTr3nde2TR9sDxE17tRHOVvgVMSm+7BxpUto5UfvV
Gk5M9TT2K++lmbGIiS8GJV3V/wgbsduGMlCswLVIDKZJGlmY/9w7IDBwZj660yh3/iqp6VJ/IKyr
Xr5DZz3wh1k3MIIcl8+9qX2TRvXLOHAmIupDrzlLMtU3VpVQ8VyI1eB1Lhtj9+xsyKU04w3g2ldh
HRM2+ulfTdmnedJs4vAoBoKM7e5tzneg/zSnJUxsL+YanL1YKBiFCyXfg5h6GpimZ3Dn/p3WRlXj
A2vyTEtSeiPwTiLjgix6IDp4WYXPhKIIUVbsBuMlugOw50WuNgcgvqC7soqv3gXDUOSOLMZvGJwY
iRsbH3k7O9nh7TCtTASoqlLQUyE6SLdIgl1hQlPcJlU4uxySRAKnvILjxmRw4kLsCe/yZJf9x4Jw
Wb/qpU3o/6BPtsR5MMUZJ2GIz+rUmXqqonCnlTzwc2+e5Vbq9npq8DYo255Azxq/cJ8ojoRyNVkl
k70qQIlsp/Z2obmcFCVQMpqMbSBHDdFz38qGynxxh45zYPyDXEIg9+2SqqpxFRgpeir+KkrIsRfb
4P5cXqBg2L5T5tjVgOeMgfdYLCHwAvnw6VhtcKti9Prwt4tdfXST25wo5gu1yQHWZwJOM9aERjfu
CMHpAndhvRtmwf6y7l1lOOpUQ7yoCmFRVrSBbTwptvXFWtrtByPKt3PFe0seteDJ64LqwFs9ElyO
MFwJD3d5qxyieje3MlyRlY3cD7Q5zUB3fDp8FcYes+ezFZnWMAUeT3Ehzn8Oy0Ouhcto/LYfwACr
JDpIalwJb3G7ZvCP/SPVRvGJzL85Yt/1d3luYoG1v/pB9QM+vGjMMTpljSs3/hUhWAXFjMgitKeb
Zu447GhRKjlnJIgjnKj1KpIwXh3MgfgJBML4jJbw4KH3kgIakpd7mjgF9KV4CKdjgP5AmVZ6IVOE
fvRnlEdz3w5i2A0iaRbaTz65EIQyD4La/TMXDdELELDqltJZbEh5sLx9lZUorqqnBioRgfQjs9sL
t0IqvH3RAnvwKAeTanoADm4WxLNYsQ9Hn+CDG6N67prYWLGk5oLY1dqQYKJeCUcOM6AZ252wMjZr
P/MAyPQUOYIsGZTWJurzmkCH+/hndapEWXGy7RQ0BPJa1EUcvH0XPJyi+0PWX88WR0//F1H92Ojz
0EKa3397G+/fl2xBiS6P8UtJoW9cZXz76bQTXRkgRDySpcH9riMlWLzzNNIkLEw0OgioAWQcvKxq
EXBNkIIGdvkwM7t68DY1YifXoCuoZZ7F15dfjhe0KGBsFPMobXRZ6mfZXpsfsxMxNUHmAvQC0CLL
3Oq2zmmALASjKx0pDQ58gUKGOWBQb8Vj5Sf7LNEbcqfX8Abrqe4pImOb/CCrRDPArEYBQIy6F3Po
gJZFZTWCV5GDKps+fQLTUDZqJHA44TRkjXXLqhugyEwj6DYuR3W2zcvUsSgpQx1DKFf+2RFH1pK/
DNt5advdwxAtcejZ3TMHdrcbgyaUejKQ59Dbh3fMpHi7CrS8tyPiuyJjqW28+dHDdyw3i3wVHnBg
qw8WgU2ucSzdhojfxVMTghtelro5YfoHYf5gAC6MpQc8rnOANHfJgsOJfnogmDWfBAK6s4tSncN8
Em5XgwgHtlJ1neNzeVO1wsz9SGo7IKWalkTmhfXc/+CG9aM55zMJqRdtoJrzMcpsLNf+bcpeMJTH
tPgvzZpt5nyozD1sSiYMnsB3i7ocZEc2bS/pS+WqVHPvRCvnUkUc2W2F20fJCSUrqSm/kmFDNY3q
H9s5C8xi2TPqg8Y3W465tspfdviSwh0Fn9HMu73aqGxsXnUdZalP47nj5Fqa4OcUibo5lPOh1RYm
uend+50fHwZQ0sZNpFyZvhjcaPyEokf/uYi1BEhcuwrMnfLG6EikZkQ4CMraCq/OLejXdXwx0Nzs
9EYS/a2XSRMTMfSyjeBHhlgGj4VWmUDWzK2rK7qW3tp3tVZCrkx+u/cY6ZNGdW4828IirjuEqjtv
31DbkSYWoeSp/7WhHNA2HatW4uYFei0Cw+a9BVX/gQtR9WGXsMP3baQE81B6ZlYzPoSCv2DT/lsu
YJwSdNEUT/jB+K4Rlvd8DLV9M4hMnGL8ykO09ztqHb2wreSujPRu897YGAfmPGwIjSDoK8mIA0v7
/2iIOzQJ9joZcRcg+OtV2b+GNUuJNmi+A02M7ATUHY+BL1u1QZEzyt/mUMGSXIQRX2aMNLNZFa/h
ev5E8zC+XTggKqUnByZ/fxDvaTp4QpQqVUiNGF2AOi659k/ywzUJ7TL2IK1jdakKZVHHAWNEwA9K
j4+vruiK3x/JShVjmoLbka/qEe4rjRU4jFqUogiWt8MUJTPXTSOuPdDBrNafp/5hgz/KNrmx3F0c
MPwvhO8u868onbVNoEf4XsTAZNdL80JW7KDPNXT2mT0QZoHeRI6hhsP79ZixZwXg7dpSEX1qY2q5
3BA+YtfqGKHgobVMb/rWo7nA6xT6aBnm3k0ZYt93KX+WMDZtyLyc4RO3hybX/m1X6FgWUT2xnOhO
Y9T287TpJtxrX8LZtH0STeVy9cFaiwJlsXO1Eo+dyGqgTy8ubWwFhdWiJM9eUeOuUlA0UhqvYRCu
nVbP5klFd0nx48bVVvgvjxhFLNdmOliFFJNt3EJygs7/Q9bEkIOhx+vnLpWA0CmPRAvAuTkVZWyh
Np/3eBUMWFxRZ+W5N4CswvtK2D5OqElS/hCcPpx0e/Zewu2mR48S+66UnffcGPSCiY0LlLPuXGC3
RcoL2POyJjg12l4qgs2Ib6MENDBrARdR/HXX/8CgFhG3A1RBVnoZKtEhGnIsEATv+SKjFWCqJaCR
BxWu/83xEf29ztlUjRsb0CkEVrjYSk+K8YJwr7LwFNLZKUufI1wFGA0zfEzQj082oiBJ9ob+QTJK
/uBZ+vUYX2dXfYX/A09dXy1fWOSSlLvjxno/dLXeZrWMTluVh+0vhfypLefiUdx1NT+N13e4fKXz
fhbuFS+mAhX7KfIbm+o9rcuqFI6NCfx06j7eHrigwup5haQ83Z9CCZYxT+hV7m3zo+seL5ssuy0Q
WdBmlhFdidjn3h2+Zu5DONKbWgjc2KuYYeyB5i1j/Wfv74rjLcgksmJn5thQ1quz1tQY5Bxri9r4
GK/J7dTKih7F5ointgQmQCAaoLdnoKdZmQYRQpNl2ainqXj/PWE9SoTgugh/N3Hh6IJP5rQgJ1os
6gddRoXhgbdbzFmghji/VEbcav7e0w4VWWs13k3WEQQ3u0k/H11OuBsNJTELbqAVjqzWxBhVBbTu
GM1mNvQWKARItqfIC6CwKKqxe129ohpPJUejRtJzmIzGMDg3oNPomokvW1Y/8Bhfub7X61fxGzhC
JS0Cc5aygK2FoE1sRmu53VAFCmYCaSbPnnhBv1atHpLxPockL9vEgOy1vQfK8OCXo3UusJZlFkbb
tLRiD2mYicGfnqXnn6vsE4PSwEcy3Ohtxi6wANiepkaAIftwMvX2gvcOQmQ/oK9XAjtccyz2vyvH
b39/mBWYDbiN0dbHMOCU4wxscQ/RwsrbRPUSfxJ6sEfvOgQxG3mL2WKAn1Ru9sF7p19ZL+y+mxRP
lRsbLBMvNQZG0+C+pjuaw/xLTKoGMqFVhTTkwsMVHOMUYNnwYLh+QSzpiVYdvPtJJE4OWmhRq2vR
iHfz67n/+5P5TEBZMud1nVmt0ieIRjfQbQR/OlCqHwbicZMckrAY2Yg+jG1bAVjySYFkxzjkEXT7
ZtdlaIdutGPsYHbOgrP0JjlD1eJUuLGSm3NBX0fxcsXtSbQyC56+XEwmZqJBHZJaQz8HlcvePoaa
rEnx32Nywwu5yJu/8AZao1uHPDZk+823ubO0xGmdIWJUoil1Ee8pIsbNVtfGslin04GI1bMjObyr
eJuxETsUR09abKW7OA729lAnSUvWob0YJdR6D/8fdgkDrRepvDAtmliCZWpPhZ15z6FshTBQk7KT
UZE8VXILw2vHJvv7HB+kLv4AMFqjduxwwSuDvVxMmye+6xFGS0OF6yisEuxVsHzxUjPvowGOjGuC
3fDUYRz8m4SpdveyhmDBV4FIsm+QrAS2/pUqOf4O99lNMPLF5WuESUMWhLWqMcZ3YlbXIgP/rxRS
FfS1+yVqdH7P/b4BNV9J3opT5MA5z24nRD1gvCu7vU2bka27jNGnr9UuxnHRjb95RXQFIQ2of6Eq
6hQg/cTwhK5XFEw/1gziWH/aJxrUKajIDSWBpdu9X7hs3PrZy1tUx2zhcyU/beHqlJ96WMvY91JZ
vV/MdFEcq7tA1O4k0BuJ9ykk05m6FVjiztpog/jodusoPVoY/Kksog82d5Y2TXVPhCfXhGzXxytG
DZcHwCQ2Uirc9+ksY97kiz1f641eLz22NglCSCiGb/vf1EcmM9HUPHTgN0K+qFFKpJ1Abe7Ep0Le
MQlUUUDhnJ4m+4Dcs2x4muGDOT/PWY2+Ux1jhx21vZwsVTq21XA/ucpAXF4Xj8LabEqaz2L7lWKM
Frnxvgcy526IYYs9UyPLRaA97H5WpkJO9PJOHbk0j6OKqhs0YfW9seNiukS/pmDtTveyhebTSfA3
WbY+SIsS2Mv4kvugOa3VGZ+10TK4+sKZk7028RbrPdebLE/lkwQ5HMsOs72fLK6Mut/a3997BOsJ
Q9x+s4wnoaJ1q4OWuqoJdRne/AASKbsytASIsHt3SUPkCn6CcT0yIqcUdnmEz/uptvMfiMndS4aY
+tFdIMHx7I9WOe2x8MM2zVJ47cQRyS+N/QSoVxeVFY2Lmd5GSPfjFPEaZoq5Nv2/Tnnbw3cp1USZ
V4qcCHvKr4ShUQoWVAIp73vFIJD0xdsNvzzG8RKSd5r3X+uJ558NH+3xwCWHpXu6y8jSqpVP6TBy
/EUtcU/+5S0c73ZUbZatgXFC/D5RDasMgZkgLl2JP41OGSg9SCxA/y+jRr1UzQ7VWZpszZluSGbk
3nvCZvBNVypkaSbKsMZw6awyyJT6LzONnMqRmu9zyZaoqzIq09Xa2UInKyfhfHLBQdk3ZbWpJ3cu
FTa5+1a5IDYDTJUpRmt9M4Wf12rq6vxxQoqHQ9EqFujGMHNGnG/xO1MJ/Sedweq/JIh6+x7ozlG0
wpXW+e1xJtUHmewhSBrm9a6ogC6TSyIS0g8HuBurP0xdgbFl5URNGVCm0XcnkHa3fol+5CiO4k8h
RVl0JBtzQTH0TxbhO/771cmEyvtrfX2DwGa00lVS5yj1jXUXfgnvuHeT0Ka3dZbnKUowcehFWFtr
Uy3xqnapg6I07idgWJTakfrkxIFup30a+P0wTcufo9HQ7jczgEM8WuQV0d1ZLACNZ5MPCWCXn8OE
BcZAi8CausXE9PCQBlZw9eLKNNdnNLHQ+JGF3A6BdDHl8EpjiqgLWDw3bPvmP08MpaUMOOx3iLkO
ovSj7i4TcLybG+Mhuf8uAviq1DsaRTivJDwoNqlD42fa96uq2g0jj0+3BuO2QVSpXQK0Q1gHMUtg
8ZmlBy8ZVXuQOEh6aAfKrTeOqFH5zVOBAM77z/3dY0CVtmUGxK8hV+LC1DJL49yZjOKqx+I+eEEJ
7A3DP6C3YdNa20mTucqd+AW5shYi5ng/P0eunFN3a+RcHGzNGmeQax6LfcECZBWSkEnje7C8FwyO
BTeMJ9rpCcOWpMkizmSweSUI8bmum+djgoll76MekD0ie8zVypqhWLbUMFN5joxbxe3yujDHbyjg
wMj6iJyQw61n2CgTJtVO9xVyiMhSyM1Bsfy99KkmRDysisLh3p//sXPsT2WocG4h9VbIMHZb/76e
YzrNcLcRbSNOiEKEbp5GoTWLwjdMtnKUO8xBJK8hLnz5q7Uc+KvMqOzYWYfi9+UNCLbux5MP4A3x
MiNKU++8PySmji8VU8wnR2x24xINdnY10Nzkyjt1LcEV+ndew8gYVStwmsrV48g+/zEYRv7eQ7vg
mAPBt7RnF9WqQJcxsz+BWOmNm8dDkjojW3ZjkzFNSjTy6b0RNi9PHVEb+TGvXiFAt1pP1pJQXWY9
GnrgGdWEjG0FRkHsi5SOcpKw0BadKVq3o+16qE7tGv7RDthzF9RtxPFGj0qkVV6uM3R58iyWG1qQ
Z2ATYRyffi54kVca4PTjV+srgNRcPYXiSTX+o7Sh7imCunZMJ3IvY4M5g5NejX2qw/1/J6eJINhH
z5HFBRt7ZpVC59qD6WUTJDbE9Wp4CFFF8bdqxp77WHnEW8yzIBEoO33TnIpakpNsHpEZUcuX+2yg
thUj69b9O3WvvoLjTMrnZna53UmDXtyfzLSSnvCddxW8I/Zsrvz2pK++oQZ1ok47W1U2Za7s7wgY
DM25WwdlDFiJoeE07GKtmhXq3nLIVLTaPnvXpStKsz1OAqmh3SzwEI/sIXL2P7qz8n0wdW9+6ELS
vXnz/cikl+6OKeuiWfmdCmwEnGxh8bntump1YgfV4D8HS0F6SGocp6Fjj5s78dXE9P5Ac/uqdXuA
HRDRrnXwptTuATv37GUPlj1xMhSsgo5UuwwmJOuzFmyvpH4w/4GYSKjGMuAV1C9bsl2fSdHruz+F
9Z4um5fY5cyx9GoB1aaCdL8p80wnlmxO796U2W4DGz7LrFcthBpVR56cS3IoFoj7S3TY4r5ZJmA0
tabosu2Us4UkcHstUHLdRjJBrjmyaZVFqD42qY338tnN8w8tKkR8nLFZJC3y0Y9YAvit5+gHzXzH
9c14NwX2VIAjYRz+rHEmvCKETFEnImdZfVdS00osdLtT6McsEu45Psyi2hS3mCj+m6tuFNmCdht8
MHdtEJTeaJVWbiFb2O6/HnIdh733iBvk8RuK/ovU59Qoa/UhVUzCQCg+eDlQNMF/6uoB2qCBSCYa
t6iU98aoE7w4ye2bdisLiIBgZqRD+LbRAqBNq+4/17hQ0/WqIZPYG+1AVQyDiSlViQfgjKAIuvwB
OqATVf8GOZVXb/J4xZbFwZWxjSeM3zIJ8hWEcFiXMGFTzudBufWZYwIe+GAyM7J5+EJcp7K3VqFb
vKTawrUU9kqPcW49rvF5nj8aPc0uGvGJXnekpqzxNcA1rf1Phy8WKtav0w/v/PzrfllkmEFpdxgg
ziCweLXw0ryn8az1wM8pQD95B/+9y8Vn7a+DAxV80HH4geeUVvAN0uauefrOrhT7vBh1efQ4Kp1e
2ZLZxIsbztNNFAkxRLEBjgB3LpcMNTtTKOBuOyI7PncGSoyNMFrP5/Aku5oyRDICsMsdrbpfUqc8
hhIkpPetXAw9enWsqBmEJiA/HxFW8pQK4Mn0H8O5+Ih9hG/K3QXGfF0G820vgOluKrz564bF8UYh
6ICv2M8usHGCKe4IKkRWieDHRqXEtAAOvI5uGOqWuP59zgOgiAcEdGCdLAvNHDmFWrNz8HXFB9xG
rUm1z9SuQyjslRJYBk+Ppp+K/pR+/uWIYVCcV7PE0ZDbf840M7LG4Uoe5vS9OU0rOeR42NiKkzs2
M+4nGfFRmRw2UuHugCLuGNGoUb/1QILmQx+PRwqx/Jq8fuu7nfjqFdmxmCkDbbqFR17M8Ko2PyLm
AM1kAS3Y+njipG/po9UavHBrWZwy1yKwqi4nZ/59195mYtFHAbsOTv5Rn1LXlVZd0W+eJdYGROyp
QANiwVupLksW/rarjyXIsmD6BFO9hZ2vx/bhVBOK8FChGOYF6e3wjv66hXApzTaSsKu8BfV9W3hG
v0KLOtapymKMNxCXLN6z88+pEvcD3b4MVZ2tAIxBIU8VcxONuCjYbzdW1LiJQX5Myg0V+LZonOgi
WHUB3IFH3rH0T48rEccmzXrDWwG/H25EnRyXTdH882T6zlL0q29B/+QbqTFLvTMQ72LuIvt1/ezl
fXoka/jr0goYaEUhFIB8oajYdjX2+eEwHI4Max/R3i5y653L7pqURMj9B5Vs1+Vi7VCd31+iAy+l
9mLzJc9dnKDsioJk4IAIM5cOU7U4VK6BKl9yOw8SNApC9UAQkwHC94h1m4QpJ/+GJz4ag0w7R36U
irRkQhKowaPBFHpWty8CJsEKUzKdYtC7IFA+U6m3ssLWamAbfeXe5CIBvtH/9nJQIZ09LwXb0Vza
kzhkeBJSuYQII+C5fVT3jMERgtJ0ruJqtJu1JRkrGtHl4DO2v6NGhkGxuzJsCYh2DhS0tRCQ6HE4
4d0Q9IOTY0v3tQwHCQuqMNTk/q70LRJhP/77sVfs9PRMZWENuLNrm5g4mILXPdMR3My3cYRyOSBN
YHc96UU3GcFeHgl6rZhELd/Kaq5TErVp7qUwbRuXrcNQDZ+6feez5u4KFNIexEhWs65vaiae8HNC
r/q/0jO0PpJpzqxaj/y9hI3Whi1ZcKQ8Fmd/L5jFKNyDCCvLXyfO4mNs1HrFPcXwpp2ICVYpLes7
7Uejgow9VfG2+KQ/0s1qFLrE/iVQJqTWIYqpy1a6Q5AXUcBdIAV0smyBLk+93vY35BMsTg3v40yH
wBx3K08AD7XLx9GUL433zYQW67iklDaBIX6TPueS7h1RFNoP0k2908tYnL5PUox0DcR0mI4ezJp6
DmiByxy/+eDm1BMCpeb8PiPIohmTa3NET4gJJTaZui0FiaVR5H4Oa0rQrK9nQwePn7zDhHwSzohe
9T+dWCVZF4YNPPjLlNAAeW2IHlK6qgCKAU17zMA7F+ZfPsRBBCoDi9X7IGZkGOI7RAAwYNJJMYZc
62S/K/Ycc7AuRkj8me6h7+asGbzvgqgGu9XB0tEvaJtjs1qpGFKkCzahKNKZ+y3LnJJyurJFU7Mz
JQ4jddQ/P3TM+nu8zazI2rr1mh6nBxg42QUXmeZ3yBY8jsRnW2hjDd2ME77FL0bBWbOMOgiwo+Dj
tC4QIiZCpYM9SW3VyV6MpIedfpy2MghzAcYlxIl3DkW6kp6h5jTPhwB0utyRYUULzVPt5G3VZINf
yzCIgbdo0XCNlGUXcntBICOwLP7F53jErMSBJk19I2C17m8K0MUqSvBLyLKRbNxcfpdbFEj80jcd
ZJfcaxXH7JI9YK+GfzdIAp1ziP1IXfoB8121h5DNByEN/TzwZM1xLpEKNLW2mBOHLJloFu1wcv6d
lWG1wgHC6cy6KwO5IqXtbTF/KW3KSO04VFb0ww3kdFiB+LdhDL0UDA1aeqZ00YY5+gfeCvygkQLy
ocmGUMpQ2AXzAfzfjU7ykF3wnZzvNPsjgxk0dv9Te+QolCQVOZP6Gv+KASo+1vns+Ttk2dpD42JW
QqDTjZs9OcSr4j9vDc9E8WNo/kSjOWmwyNBWqT24C+ABX4Zof8Ip6Y8jT0gMXjM0yAaCJZj1R/DM
rQGycju1IzKnRWvYXxsTbIYqZzaNEc9M7T4xx2uZjhgpP6EgggyW2+RdICmdEYX4bZB/n+OM3Hdf
L8jCbxApxRw8w5Lh6vLUHS+1BistIVh0suq7NBncJ6SE1GTiDQowUz73rF7+JnkjVz3Dx6ldRvs/
ebxG3LPSj1onz5vEIqlcuPfS4bdpC3q4sE6UdZci3leTybsroX3NBWG7x6MY0JEVRIxCV5DfF2Ew
LeO/AaLtiITxITXn0Uepoh2WJ9bLoD7AxdemjzCWf8CAKDNpEy02nNxYAWElric1dK8YBlE/7kJc
mEH5J7u673SEadJKZJcO41+fPysXnoOnwCvtA7RCY7jXj1iZsCDiSG8SXBgrgyBSw+u65rkuWTmk
r8KOYQlL1hq2bvjtBN3ATUtd1w6P+k9Po42ef3ri5KD7FzSxIM0hnI3GgA71gzPDYddS+yEIQ67O
LMNlSSzibBLsow6kg1eHjN0faxe+2QS7IAyGCX4mRNoYmaYBZQt3BsU+2Hr614cNG2dMvtxeRcto
Hv49l4vSuR//afeJGxSBNECzm0G/vOLg1KjvswfDIydNnEwyj5bEtDNXShDjaN6zZ5aVQpUBOCJe
juA+47Tmnf1lnQn7R7lepX519GXiZcYk4ieyoUkmtji/5GhzLsuqM556gAofd0ZkaLvREWcvSvJ7
il4qQoDZz2GF3FEOR2ivqJK2JONna0eDvQTrvM7JrCoJzTqBb6iwPGEY95NkRO20tgGpORs3xjBW
8G8LCyDXoVSlE8KRHLowBdRWPwTfaJr53nEoD7Ze8j4aenMVGTGy9AwASndfhbUDWRhgCLCnbqns
nQHNReBb+iliwNa1A2ekPUEKHMducRDHSpoxs/RtkiyaS8UVxWlkmRNQ5dfIUXdk6DqYY1KWbF7E
XtnZE7jjP7SAw3ZqWisL89C7uOtANH2Wa8Vu7RhFBCYzSAPPh09qT1oTNP8UYm6Pv3x1CZZaqO3J
ZkMnhF484Q3t62kBHvH9PcvY1XeDyRLtxB7Yh/1SuXLSQDtsHXcWPgQvpf2N1xz6y98EVY9Zv+8H
ms/AJuDCLRh0K1XtupllVQcvLeIwVruSpapIhxIBkpIcbMBvzb7LuupaIcrigDDiNe2gc3D231si
lc74fauHWcP4zGIm/YNq0X63QjjgU0wDOt68659Z7eocLbFJcUrw9gYIsrXvInteaGLww2LIVcOi
sInbuhU9V9BNzF7G0yYpYfRAaHQPXwTv57nXtM36qosj8DlUn+xk/hs3ofeOXBghsikCdYhmhR/u
/ZNtVuqaVPmrzYzbqTl+6dkfNwMxgPYF/rka2b+NeLsgTlYpOSg/XBEpWVAl1oECox9wMxLVuHLM
RJ+XLZIfnPJ5FjRHVxd9ExEa2gOFZJEvlAXpNQNapbV8/Z0XI8M3JdoAND3zcTLUU8bv3GOdByHG
/rjiBwk27uy2f/ENpZ9H921/oB6Kfgp7FF5g6sqWaH3YCBrmMhN1A7/sFOI9PFp7HUgWjjgcJzPW
diw0HQhq1GpUEN5gLepww0gAaOD5PKDLHGBofRWMF8xG29nqeDpl3WHRyjxlavAgxcC0n9LippFI
TXiuSyTN+rjKj/u2B982BTQgBJgdwtV11SkDozqfYHsKFMXk851HS6fsCEIZlikqzvtVdyZ8B6s0
PJhGCV1eDrhpTjvZ8TPxdeaYfruYgWjOg+sGpFCOqJYb4UzA5IOvVuN//SJgsScRvUqeBUAVxadG
oneNI1C5n4yjbFKAHHD90ZUlhVBSUDtDm/U01fPrZeSkDO0AD/Aywr6SUCdTjIKyvjg16KPleWl5
+62uQe7kqTmbuUnQsiBavqzPJZVcgSy0+EzBwBkfknRNWXAlwjDHNM7KBNGigvADqsTBm9yisXl8
xL/oaWsjqh6ED7MYd61p0fGfpLHOEjiXBDB7/QD4BbD8jIJpGPF3eZyhA2vcp4h2f2On7DhLRW88
bch8wBkoKlcCdBEzzh2aWdL2WUfNHdYnmnnzzq5OOR+YLxVisuhJlFXamwdsudvV9PWurM1AmL5b
O/O5Ycm9uAlYWTJkwNswaI4ZitIOhSfX5KNYR+OzxMQSTKUdhDHAfh0Sa9ggwP7+n2nTeci3ZpQI
c6QzKW29jOkTC0qjLDGg8MDF2a2C+r5x/wUFUY6Onsk2zxdsSGjU9MjiAsyiOCKUOZjrbqgxCyP4
jxhvKkt8yWo7pk9tZ/ywMsqukJwo4TuKgQmqRQq+lKuds8Pvr3l915t1o68naMlQAb5mlHTx7f4b
nwwASPzBjM1seA0FIU/KChdnFMWvb53btH4BY+8B8F3BCcepBD5/ECd+prRTeruaYNQr7svzZrMU
LuuWDccsWFs0APRqyjiFxuNXsepWRBi1S9cAy0z0b02sc2/HovVMc8RySM9VzrVHg0IZiS3EUIvA
UBMdGjLNJm9HPTx3Olk3P5swq5VFSkl42GMzpWj7YRLVMjLwVWUhzrc/EW/uqicazQJqKyxtlAgN
+MZSent81rR4PqRS3NEqA/C9VGx+nj/vUMZXzqjMxA79yJfQHss5BRsAVpT52D1lmMpanKy4VJIV
WaVUs7kSf+GZVFlPoWDIihU0siug81XJWN3imnG1+exomu8GHAlv8U48R0YYbfDlORD1FehDCs4v
qX9RH3Q6UCmtv6XvQSjJ470Wqmb8eZQGipTlZ4pKFnKqkyN+evTlenUP4oSzBIfgEctQhdXz48Bj
cCEoM6wZYFKsJbERWREQ//TIQ2+Xtu262Tlz8zS1mWngiojum2m+DDhcbKNZEplt1CuLElC9yWTw
kvSzf/JEfM0hQm29FjllHnzE1mRCuBPYlBlTbwqS/iEeHC1e4msHyM9cpM+b8MAae01gl6uC6FD0
NcSMZ91gkmmSDr7tAELqTXsag4CpAZNbU/Tck97Y9NTclAHyrv1pBzS64El9kfKUua+iboUjYvVR
0mxDzC/qGFojP63b1ZXSHAfogXSDRfpdiO3AX8yarQVfHdiaaTAz7I8VjXnYCsOjmImU0Q5HY0/q
FB3kAd30oGFk/R7fYiDeppw9J1PU0xzWBmS5mZYOlEzbHn6v2IZ9SJZbwVqQKFwy4Y6QmzOb6EJl
0B/o5lNZ3jyTT9D6p7GYF7sWpbh0TyAh5knnCDFrsZpGZRHoBeKlmDwoIALkkgtIwoQPbQaO0Clj
dS5hJiVH8+ufiB96RtwUo0ZxksVtUI+XTxoCbJ9qWo/45ykpaqqEK1OnNmGl+uMKfcKlYJL2ciXH
zl5udbqEDxu0ejaNjPvIi3uNl61xYG+XjvaQcxLjYScCTlGU9bLMH6Kh354pjSWqzgwholPjhJsO
qnRobHBmtB6DfpZdrYWgh/Fe7NRnXFPDQr/9PbNAJPy04Ll1GXiiSponG3QrmlcpBkWiuQMC62zE
1Ddzi/5LYmT/dvQwU/Hw1Eau3tU50A8ggbI/1mC/h0MB2q49q6k8gu34dAoZOPcUcZ+am39nr6/g
Q+1+WmWbw11vPf05Te/9emeklZXzw/65m3a3YN7HGvzaD2gZ+7Xf5dK1PvLNVVSp6IA2TPTO6h4i
6bQ5sbjLDjRGKdkqETdkqs591wl7Jcxr5vLLCnu5bH7caZSc0+ELoM41VapRMiuerX1BYvc/QxSS
t6jffnMhaBgZzcdlv6y1S4eVPrSUHSAk201DZlKfaa4T9T4u1+vQ6/rnWCpn/7rLqNClgT/ucj35
utZNglGLmk/j3OJdynRkNHa3VHNQS5YUH7OHdnn3NZ3cc0AVLSpHqYvUIKRxmaTJqHcHj27Fsx6g
Aus1hnrlMfKT1lGVN+gM1q6irwMenLr9pG5bZHVqc3KidHhWgawbNoqyMWEYkWVPSQIGhBRzU3BV
eVBTGirVMgEd7oFTZ26vVzPe2A0C9l/TfutbzEhipmIUCu85DANyuhXAZT/BiyVGpnpMDm9O7HO0
5TLcP8f4u1vyTOCVdHl8Lea6NdEkTG6eW91FQNZFaD/6lxJFws2CD9gwNYuSphta8ka7qYAVrkXk
lNr4i/uLD3hYLXBvfdSKBRtXyKtvTzms8Dw28SvSYbnQuQ6R/5uPxuaxNaypd0VXyrzYInbydZ5P
XLfYhoAJx5IQ4l5QXC0xs1E5zoJLAC3noBo3LUSC+CMUDIWIB/441NtvMpKfLQXnyeBKUW8pchnY
nl+Wi1ZnDoy9p9ot3Fuq4MsUJ2cNEGVi0hcLZ89HHaOCdO/HdUdtJ7P3BdLcd0ATV9PilqgKRFGH
8TnzUtZmvVPCbv+jaAtZMvVfn4bRKxqSM3JLg+P6JpjcorpQJ/qV5mxUvopqgmDmlHMoMH4IsjyD
S3c4WVVCyJwaWOHM9KZbMTz/0zxBgI6qho1kK5+8luGWIE8qvnn7GF5v2YWj4AS3qxBFpJVIYUES
yWkYeYBpspiD10J+bctZ1qpRgszgTbSBD448PWGlx+uB8GrXhl+0GikazYhYmrfFB3PBYC6wLXpB
jxDvE403cP4yplGbmK5JK4sB9/ZH8rqx//EfEWBhp2UVYXYtrHOGd9LWEe0QpjqIMQq31FsXZPCQ
ekCa43X0y087aQt775WULiJuaf2KPT2TtdULgRoFk92SXd5jn5eS9tjOHgyaLuiWsyoI7NTEN9/8
UfGraLAvbVspsMr+7JWQilYP0UR+hrCKkwG0n8K4LSLTmti89aTKFJ7x3yXp+T3rzeHB57FDCtiF
uFdP2q6/Gv0AVPh/rDjR9xIAkzSxwlb5stwgd7QzlXRG1uyIoDJtufioO+lBF338Huiz4X2t3m8L
XSk7msVWjfF1q1aAC48l0/ScX/6nCiPo/yjCREB0zFqeV/+FYZZs1E+dBOY781KeH7h7ua99TXVJ
3omRep04G44DXZWIPaMx+vKxm8jZ+t7TXKaTT9mUdb7BxC1c/j572XZl8/WnXyHM/Ne55UQr/fqR
hXOcKKFyGK/gqpbczKOenjcKhOGj5cNQBkv4a9vYSFFrw1KutmUw1l4OonFsYQqMf7PVqhMwZ+jG
BIdObpBF6ateFFXPOCFXnpEF+5wPlqD/0yxFv0FGh5eoCJN2kOd4VUjjVAdMVYWLhq8lBijxT9Hf
p1hiKioS548ZvCNk4JGd3/FkmZz0oLGdbztglEgZphFth+Yr78v9JKJ+wcpd1dy8hs7QRXYxH689
YPrI5yPhRxRGM+VpCd0nNOYP/nNAJ2gVoMLwi2e7lC22NJYxxcGpv9IlKIKG8AteeOrz2TUYje99
D7L20Gd63LTGgqA1ye0Mvdkyi2wQYgpEjC2UFhJhI/1mtVWN/YSnh/LRMhB24pQ4eyL32S2GcyRG
vI6nKxM23hwMKytSygs4o9Kn35oWmawrhS6a6if8GD0Kqeq5+6xCYsgdMnE7pNmkryVBmt8Ce4ac
cYJCB99gbWGFtS4kyMUJDSrmvgIoxbM7HNucRuOoX6uE+SJH7VbVbdSj6xzPNpvPxQNhGKkKNDY+
8RNnQWwAUzDOpxdivRZ+YavxhDEWsyVz5BFpDmdbuFi8AFf5hbsSTRJ0eA9Bo48hAo7TUF7iYry2
rDcsrY6Eh1Rbpo5RFiSsk5zPn3qp5EdMWUoIA6GJuPIKQp3m4ZNQjoKiiXtS65hz3nJK+VHvwf35
PuaCe84+BbJz9LVPm4cEEIbS8h9mZH0rRHF79LlfocO/xcKQDvD3I87dGRzpgNo+RhBEuR6ffkXi
gUc1dvTtrWlfZ63O1HFTB4dgFGj2487tweGi/1QmLURpFXvBR6iNyf0/N13dMrcM4Tx3fERBucqv
tilRGmSV7+m5OVy+cA+OCAVhQRzALEHpob49FLyvosRSzmkzgPkAFg3lCw4TyAgWE1iaXRkvURuA
5OgKM2zJ0Czy7jpkpmJr2cnXoO7Yl/iLFDCM0barxbDXzpvcuwx5xQ9FTlz2O8wAmJJ3u/i0PvTH
+jTRSdY8bBC10WfwD8JhA8qe2G83ewRfT2w+6RDgXDpMajriZoC+HD+q2UoMg9zYYN6DTZzeLNT8
e9PEWFW3VwDE76lm7Rbl5yV8wA8a+BXs+zyJ9/ORADoO4p3AwJDNYyp4iQkRT7cqhjsrO2TVVLsE
ruOLWoRjsZmKc/neBak+dim8vtKkfbxpVI8ub31ikRkIdAcRtq6gbF1ynKOwDdcbV+p7vf/+CcS4
bztiwOD+Yt3afv3EzsP4gpfBUHTPTwLNiNqIAy/qMIuhksexDD8Zbm/jYyhcKGkarqJH3p2tjkkU
Tn9RjmOip/BqmFSiUsMdSgldL1zf0+CqAz2VdE4FufI7SR8KF43ywlIQ6GSx2Oo7aKIOkI3XBjZ8
+ion2J4NB2GPE8ZvSKfxyxfZpoFP3QQ3vVrhPg+2jlKz3CNWucNNHN4vneknwLisJKqoIQ7mBLIL
0GI8/ihETONAaZyCZzK20jpMxeGwi9hpLbFcRTYthUUahDFH78qBAVjtAXRDEfPjwXWhg0tuDssV
WiRkJ4T337tZ6nZRToQFaBJvL881mG9Hc7kiNlnfvY7MjwO6Spr36fJUHrrim9AkERUJVpesbTiU
VHyOX4WSLeP8UEGvRiFsy87Ulw8/TVm47s2KjEWtkOZ1Nwax4BX0x29szfOAI6tL1AHufiDOMx7H
H2W5OQgdoDqlcUYGD6LV4br/Qp/CdB5HCVUO1Hk9Z+9/yTiMiSyc/8bfHjCeMHGZWa3rz+1PtHMP
PdXSy2mkdOo2GiAtUvpHfkvKjLyRqYa9Seaw79N4lzTX9s8I9Dn3IpRCrQplzAuJf49xpfb9QtkW
tIKV20qoANAeY+q4L5RIYDfvj0BAX4UST9dimU7K+Seqmpag5FgrXK3DlnRg4RBtj9y4/v5SXXWm
Fe+XYleDnboHDA94Qoq4FSdHKFUKLMubOrSFDrikk1CHtRDtrw/h2187k49fYQKxbS0guR494Eo/
eDq7d7aGdbY+eUm5OYvryRJ/upErAr7IaZLtLxU1RwZByGmkcCAxfovUVcKQN6YWp+2DO//k6JSn
+RX3D41rww7G1k/ZxmOlh7Tn4ayUzC+iKB2VSqxtIYAtu1BiVA6LSEQRsFjG6C9m98J29i6FvHd2
OC+wRqxr3EwNm2FJzIAcSApL+8HXLqjs1u+qtstABbXx1+9+VVOSg1jCT+MNzWL2ocL6I0cWlwOI
glVdACfJ0cE/8TxVfJ0+NV1ebLzYeLX1cpqa/13R9kCHGn6EnMylbU83KK6T91+U/iS/O4xERWFe
CVV5ddzR0a+CM+zR4EeNPoUFwvJBbz7EDyFfh9Iv/wQFbrQmjlkE/F+bM+jwwGTkqEUO5ogujaFy
kUofVhTgH7yfte0nd6llSQIs+MbPyBM8NAOjUq5hAJieS10TK9jiQYd1ISJ7q8uQkHw1hsIqmPuN
lquBPX33rps+hIwYY5bW2lV5A6Bafyf6Fh00m9jXCLNosNaRnU2sxdHMeVVzo9I3BHMRa1TadKOQ
QLe8ywCD0eLQSZFB/t3waPq/7Mr6wAwsdEcSkLkJp5BcQxpNneVtXah3tzpyXHzEomjsnL0DToLF
iA10uDqlRsUCc6S4+ujfdcs61XIUErujG4ykW9JLovfwKYNO1jHcT+ZGadBDZvfWBMrcW+0ULIIp
AkuKmlG4nw+1KM3aPv5qbz7DHXUDi344aik44i90HcbXQeGFf3JQaEoTJSdedK0nHLr1kdF64wBQ
hUxkmmNOzq9b1stVKaRb5iLHEi7nWciwOWvape2UANx2plqZR04VgHBtUxKbW2+77sp9WHoZgnW4
4/tXgRp3Jp+WNmylF9x7Hdukw93QjqYDW6nsVSi/C1xarqePc9NBq5pzEwd/850tXeyEL0RqDvBF
MDaQZzNy+VBejfTwFziJxnoXpJrtGBteVMN3zjlX3s5gMvlEc01r1jr02a1F4yDi61dIopyTyhY+
mgTLmg7e8E+fZjvoQrm8En1hXUphmXT4Tziz4+PcZfA9W+a++FvtcTJNBFSlgIe+k6WkbpR3UUD/
po5Dt8yyHXdaNO7nktzuHVF3cfY6c9OKWSQIp793je+WyM9yC03RrxcC85ZxbwELNqC/el+vnGDu
zT0O+/soM2wWM6a1tdZf9LL+tu+srDlawFCVyYOPV93pU/UEVJKwuh71mWmrN6CP4FDCs8ArOhdI
SyC6DIM0bBA7NE5d4aeHMU69JU316Rm8j79MgAXGGiPRUaC8xg8fX09/s4DrOTCNenFIphIol5/l
t7/VnaU7geygGjPQ26xbcERn1nlx05wUWotec3PVunwfg9rRMHfdYM6g8bjtQW/BPWsOiihtQYzg
GjxfdFBOHRdnOBEh3ZtOPtIdnNOsnwzfcB6a1QOTrmEyvlSbgfK92nZsetSfeqdnmk/1RAQfcZAi
3otUez9Tg6DhS3shY8PEa57DqssG8Hmuu7OMPZNMGq+c2o4ei+lEC9NHXH2J04i9/szpE/gyERHi
9qIKhG8IJ+KWUUqtzrGb8G3X16wtqPTmwWLDKZgUCvxHJihCyQwvK7UQnKwoLXPJBSohK6u+89MY
R0N5ZSsFIy3QVF2IbeSCA55/b36QWu/Lf5RgyTwXZ6sAWCcQiiBPDt9bH/OSMskDj6wkbsw/ErdP
YBj3Vc654HiAoTCQWWGxYY3g4Lhxn9GE3Na64u1f3yLHv+4I5bQowqYJhqDSOejn56kkFqRhOMDk
+Da91EVNFRv3v79Co8nbPX39me8HgFOw39iIzxsMLw8M4AQAnE2dNDSPSN0+IvZ9rI8L4G74l19Z
oOv+FV5AhIlsU2J9zJqKgAlPFtVHSbSfD/5n5cHZMS+EYAHL5aZqe66QcsmSMNEe0dQy8Vv/DQds
pI0ySbHR78T/ps3+SpjtdESVkPCVU6X+maFYgLjOpMRZ4Hky/1WdIEaNWUuG8S2B9/xpCUdwe/gW
vHk5RWXQhsEH2eCivYCbTjUiLGFb9VzoPd/ZOl9KZBCwqtO5qAipkeQ/Z8rAw0srpV7HbyMC+8TG
Yps64Q5t7aTuDYMi4WFjhjbAiD0QPpUA/Bfz+q2X6lrykE7MNUoMvnM35gx+Tl7UmbRiqo4i9VSp
LoauHH2QdSnDXhfiq7xe4mEDOo+RWHcj/WFxjyTBdEYT09fUo3u056SfRvPBf0uUessLNulzVxRe
5ESllNLkV0PVB7CDJ5TaqMUt1abMyIDqQJ5wxk1MrXjho7Xa2AENQRa1lLk19+IIFfU0245pLd3y
87k8DeEBF+xSzkqBSrD0ZkCIVV2+yflkgnE78IUPWJv58in3D3ar2WWWBf1PuuStl05n8ARzIVpX
nzX2t17AeJhwv8TurIHlDgDVxXdSlQ3uUiZki2LO6BDtBhF+2Z5DdibZkoAhgwhD/Y3wISmRWtRu
0/HYjeXLFHH/YSSjzRU/U+PujYYhEstC1ej333zXA6VNhzTTnyiTk04+K8tC6cjfpyXkx7pG7YtD
veC5kNDQvnURYNFGIsDkZtUcEjkOJfq4Qbx5IVji6xwJcoRZOK7CmJvr6J50ktsSsLwY2ATMKKmJ
vsIqNvnAQ03ZrGHAgsRmG7uS3mebdY5IwW3hERxr3N4nx+NOqv2hkza3FwfYp/MkEDHM3vsNyYtF
eHOkRcgUEokZMDME8j2/dweJ/ozqLOGzGX0xA18XWu/V7W+peSF+bq2UOI/xV7Kp9pmA0HDi3U5d
01IIClbe6ZGWtnm1O7n0lY5zSx1vW1kNKgUnsWLqaOdxvK7frJUKxCyMb571ywVsdhPBwPdD2tMS
5g/LaNRRUS1uL10FfsrPm5xxUIQPzH365jO/ugiXmyV1+fba/PlpdXKgBxyE2cJP1n0Tdbqj+MtM
zxbfBsB3WOVApHQd5tiXy5JspatgCZGsvDHOvqefPBazEOdGclCqNW0skYRc5rZJ6UVSb0FQKMhL
IYl7tt9vRj42rHcsc2WkUYcQuGZtJyK8q0Dq2ouyq4zLwqlJSRVQiemBG+FamhvR2dAQNgruPxE4
D4Qio6sVEb4Z+mDmyJ5twZcvDLhd7HKBHXMUsPuzoZOXNwUM0jol8PxU0HyIKi/ZxDqlzkuBnhOp
Jg3QKQ3y1tLfjurleHDUVrqcaZl1KuSDnbCLDta/Wfky3ig3+idPApkocNDDtCI1jvhDaTgSYqub
B+3SrkQfqAtD0Ly3bbfijZfMIFbGUpaDZzSnW8ZS3ePnSPXOf7dYCg8bIGFg59G9cqXwYCFTsGg+
0T+Hq425wRlktSUQV8XdTRYT7c6NPN2vx2Mqq4+cELRsqMa3WtvwHvoEf3+dorsqZLesS75meI+y
9otcDM15o2gqcpU6OePFD6ONagPoeEBz8QupfeEtCGEZzJQmqFcDRzjsPnqSum6+AX7VThxvebV5
nxbfgoikloX7P/nX/ZTy/w8oX3M8gXG2Te9YWTpBWtyFdWgh2tKSNo9dsSHMdB+mH3PMcTqvF4oU
m1huuzihA06wHs+wJpwDXh7xs6MdnZICbQZUn911qSwqTzYOkuAArS63eBjJ/pz7HLjhLTaXLpBR
eIVhVOcMhLBmDjv2kpN5sDR9df6Xz42ZVBx9gI62U2EVQmxnanJ4ruBpkkFvmrBqCUahhs13kJEZ
kSXJrEzF2oI3h7LoVuujryz/RVyVEGipiyuTxbxbfgC/GJIDrg8IBW/Ku0jkj3H2P/EogodoJ9+z
0r9Uv++uQpaeAQSAui8DL61CoGrz7jBqkTpbnL/ubDMtnIFu9cShoyMCtsf7ONMjbiTAnVr59IfV
l6DxVap3vG6ZAgS47E7p17ckvn43zvpq71gi6I3+0qwjAFdAnwsXKbmlS/ywH9aHXsptUYF441MI
FoDRtF+FRwgZU0j+PRv8JahssmVc6J1UYLknm/n5hc8752mfYrHcVCHLqQSfJdF3tCBXbI2WOeOD
j1FVDlmddLrSu8gFv5/w3I5lW2gbBFE+/WqEaSpaqHBYkK4DevJPX7cihN1n27ucbIpfosHxd8OD
TLiaG262kpg0yeqWE7rhc/hHpdJtTNGbjEQf0f1wZ6VKf9GRmzsUtI7emXMagtbIKDBLZd5C46/J
TXPuuFPO9lztqNjDnk24aJ3LkvXcl/eD+su5MvmSBz8sKqpyA8rtJ4GlBlEtcQuga58lt1S9YzyD
cg/ij1vijbNFdoHMgJV21aO9mv/GthYJ0dTDmLwu1nDwgN2Kkn/O3tCeou/9hTu8DA+DkibGrJR5
qc+QwmMosVsCNAWyd1e6f7nEHcfj5Npf+6/vAkon32Y9TfxmwNy1/C73WSKDvugBuVbIWs9SWVIj
hArr1xr5MIS8BuwS+9JT/komvFE+y30emeDpDNUXzE62fBbTGcDLT79zdPT/9O3uJJJ5HJZMMb+b
Rs7OsDy99tHjHk6+qzGueT0Z+6pQxpRA0uljyjNLzeqVjIk7+xbUeoESeTbfC8aa0lZGISts41et
ztf1VqJyKelLlY/IVK3+dUfUo4PgWqeiVzM2QPVxbcHeV6qDJECp87nZx/IlvN3FRDBjBx8dzUrq
QdKMZN+HPliJ6tFMLcQJ1/QkkU0oM7dVTM2UtL7q/5TBqWIXwJSL+IgiCtkt9WpWqpPaioXlHQNS
WRH1jKsWyPk14Mgz2ffUPw1FqDlCVle3jDGAdpGanT+RDm4PMGQur/Cu6LYy9cHgSN0u+dggRWJ5
+ndXAeM36/Nasgh445bP8HxBEU9KMPghkdPwAcg5AAeS+oXZ8y36a6HvNVZJmIWBCFoz6iG+QIRh
0YdQcGQUMCQuu8mlWlhxtXCHanDL/4hQCTwN/6713SMBXuVhUWaoP/I0NhM8VcBE4Idh986CZym7
C1uAi6+TbRhZor4sKZ/pGM14G72VWcms/001t5Rs85mbmA0t//4yKqJ3VYMaP2IrZlfhRUAX8qJG
gyxBbmPDODD4+8D2SXIulubl0cMELDzWYWQ/Nl8de0vMuiwi/AxDnovHKYhj8QYXCteKNZVYGPpL
ObsbQ1IYYOAEzzbVxLzYVUdFBAq3OFOxNGkee2YsB8235vS+H65ltQQUsbw0Fs4RbiVJeqg47ekX
9zm9bpKjh13PUrH5WOwF6XhBEikDkc3RRvzdk7EKr7KE3h9dT9Q3ViqBsmbAQv2TmjYTjhOyaI5b
PqntwFDNDOJLUyTd923hcLM/d5bxoIWkkAOB532oQW4MZtw9+58HXA7mlh52+R/Iy9SzXk8cnluC
nJ4aL2LNVES6ae5MGgKQY9ekxxtNbHS9UpmH4iPIDBiJo4skkj6Avpqfii+hO5HZ9rSH6B37TuK5
tx7UquiwbPHYs/WA8HQGGSF46lhcXfhvMasjPy3gN3zh6qvX3umJvrMqlXeaQhPuiC8Zo6eHWTRv
pjtaAJXOc3A1iQ6yFURyBuWFkiHTQcUHZzbtEVSqQU0DwJQPxKgMn9k5aHB1qnTN51OAFqspGIrL
+L2ZPsSKA39m7aoZiZ6kB3VQNF7jiQ5sa5ewPd4nzLXemhjyVhVSRzSxoKDcjvUT5LX6gm4DmXqD
cqACs2Y7/Bs5a3158S091GDk4s8ww7umjgE2X256F+aITUbATasHlYo7zpLzvD+erif26ki3/4Gj
pQKHDf6u5TSUjk30P6Aoi0IP1i2RniQAfNv6CxPh1MT+DCY/w1Zb3t5Q4MVwV6NAljPZJlGMFKSL
uUm0w6bDXaodxnvgDI2Gdq+Exgx81z7LayMHfgN1OGqsmKG9iAfy1qlVWey954bV5hR4+iHKnovB
k6rEscTzfqTk079RW3BpZVgHmC+HwH6cETpUKDFYjb+wDB03+k5As/6vlJ2/tJzUC69q5zkFETHR
7vbPzuncdy9pA/aDyWurfLOgR3CG3czj3w6Y0oOF5k4QEYUmZcuCjmdw/6o7m373Gd7jmiskkrCf
TgCWkEFI0+BN8uDVFrVrN/obebU+8FsdSpxXhjpZnlvvUHa+NxJgxxbDcAy7bU6aiK4TLhBQMCwc
U89J4aMhU0Z5GcR2aYMifcaqpc0Ygdy/VeypCChyY1uOsdcLtEJgwRukEudAfiEc0EskrfSD8hgX
0EDXADNR1yIS/V1I01ycRZhN6MEvZ2c37Tfmq9g2+2Hofsma85ejpIcj9WRzpDjlDcRvqrWY1YVP
0PAZSTwFqfARzW/2Hp7BRnyw7CF9ufVTNo1JkdR2v2TB7fFe3FQGXfnCTlQ3pmODJVqcm+mlbVpe
psQMQlpV3sZEuCX22uvcWAy3EZj7EficWjw5RyvOemiMWs7MwkCxiweCMrkAKb3CaF2f48e8vSWq
lmPvsxTmZjtZTEJ23P40beK5IhXymgrvxc5TMlkV3V3NTzok8goSRI9C6wz0PW6WxPnVDZHiuPE7
tb9OSi7beylB6dtaXK/FPHNH3qTcGQ6KTIHZjLsziXLyykd0oxaTC+GaQn37IP76SD5PzSm1b8n9
3Pnf/vD2pcUCYs9nl9Afuit6whLKHUu9dlN7rz+yl9GiMnGr0OkMtPzI/zTv0v3su3LRjY/XQWea
rm5RRCLr4FjVxhBxEmH0RBNP/3E3j3BaGz6McrExwG8B5kbS9V2oiRHHv/NlKwmILsJvoEQJj8Rf
Znn5NgjsXG3rLiBwJPwk2VyBXGqqBgld2aKYC6YsAeyN+JQ2ZtdjGWH5Af8SkCoeXegRfqw4Ue+V
Lui2xbQnIswxiiZbAhBAscrQdhuVuj+FlMGV1HK8w6DuQt9QE1itgOT5u/ruA70BR/ftm2vTbD7u
yZ7EH6g3QRg2jIpHhnCplCkMuW+1wiAdFSsvqgqqLfxlDS4LKbcWqj31SGKgJu6f2gOCJOWuHsEl
sOCXeySEG5RT1E4FdAZpBljyisZ9dcTRgfDOdQtOsWsAm9OKeSvZ5EPb1VmMLiGiH1AtOpWVywEi
xMJNenbIhAjB9fcE+6O126PWf751vOj9rzMfDpjOLmoe0KXfQYUsgocKWftYi9sWhClt56yPbOWz
yOhj3rGUPIOO2SD54AVI4BO7uC+AN6SYsiS0UWd+xF9CitMQwNDyfwjf+6dQccAg1VxOmYgVH1dk
AmCVi7+LrgJJbeMJ6Db477ZUNuEm0WXr9H4jo1+IoA6AYdkmbWS+IBS3Bb9AMn7jk7q69WpCsocu
RL3uzknAosXHFS6fjRV8YufytWfw5yeRPuxUCCZrYMmswbyPTLdkNGjCYx4ojFUq3EUGlj2dkwN8
Pt9G5BXL+WgjmUKDc+YDklYCb8jiBE5J+eUBs5qHgaqxnqMuC8uNxrcVS4l8vD49jMlkjVnTV/7R
Ti4URE9SbwjisGzaCiDhFQR5OZqvXpVw6qsqyXhQpuLRb+A1uNICMQBUnrambN3I3wt1MAvXcoAZ
8ApbW22SiGiBRpY/g4kIHTAy6iAeVF5T4biMwkU9dfAt7lu21oAZeqpdN39Rsjfzniw7Xi4tu+N2
0FENcaahDhJnTTRqEHbeCTJVON4vujJP+8P4KD1jRMGoTBHGEH/dSlf1hFSiSTANjFaWiquYIEgh
EoiJ8NYLJo4DTE6R3N+BxxEMtUdB/p6iPSMmZRi+4EtAH8qaijNaE8TDZBWeKx2SXyiZdi9wIgu9
qZLg2Dx4XcX0rdZluzUNi1FwvC5g3xfh1D3uuDKvT8bgvAAxu2cYnXTDcAaXcg71ahkr56ZDCmJQ
mRbDNGFK7IyiZLZdCbyiQMRJpzjdIXDgfHl7X9Ic5EiGWfz+k2FfN5Fp4d5h159DNjIlSZjAbZyN
bliwDi40+lBzb9o6ii86aRor5LaFa0Agx7e6ZR3FG9ScsoGF/+nZlF9bGMIL2OxbL1nO/P2POg4u
oQOKq22rKl0PBQrvJ2IVkYOoWRhnaxWCfCVeaeLC/HpzDRFml4hdrRn9EuNRYAWsCMrIqGZqKbYx
9cbZrtvBvwsRcZgeXh/FsQIHQRB2PPnKOVve8wNyIX0Tcx7qiIBcZen6HZKCWA5WVs4jfDEJpFW3
MDxoXUsQBEhwu4PjA+hnH0IasRXZwnhqO9uXk76KLpzkjHcLn8z2OVvhRdH9pmM2dYLTL/YANRok
PKoeKuqnL+5hKdWLng1DFEOPKHxETwm11MEUZCXw7HCkau8eTvY13SqtCwKtSzoZRLWreOVBJpzG
T0DN4cqBChcDelVBzS9o8Qv4GJgqVasptLPaYQPOd3H919q3+6NP2uc1+KJryRBuMspD6kb1enT4
RWzskmp8lYjsB2KGTfecljl9nt16TTk86WSaSO2A73ltqqwmDMFoF7KCcyK2NnYG+K08EnL0eZUn
vwMeIju6m+nFvSgPDYbXEZ6H+CTCVLtxbyjnq/jCeRDxboqPFX3BCBId7swSc/HPyWP+KcaVB2sG
JccPgXBf8fcaRo4iYUop6hlOVjBWbxm1NniHE0jjacKYzdnJnX4ApKm+6A+YXz6fDS/DwgaCLLIC
d0pS6UsjggYwvob2A+nFxqT6ScxfV/G8urechnJaBhnOeHcvil8nxGDWBFCJjt42y2R3DssNSmWO
773QVRsUqlvyFF83ari8Zj0b49mmO34e4vVQXjD4Nrvcaf/kBSXUnpwHYQstfSTe831PpUNGQoHo
PwtpIgc6e0ctyhh7YJ6/2YGCHTBjOb3HpnsrVvD/x7uYz/N/aPvSaC96nijuGFxJpnLc9UOeY0RK
nsrfOi/s9KUqo+uLGYqE2bsn+75dclfeTIC/hkBACpi+LvZ+G9rs16I4M4Kndx+6/mbMBSjwHj5k
g9Bmlqd8C927EvRCp7wgLrOhbzuDCWE1zwVtXxpD6ZxXyN65itX2XIjzrhY9gAG1XW5xgb7Dud7x
prFNS54R446g3NDrXERfLjdoWbq2ih7GLUIaIEYWJsQ5ETiiV71PF4w7HWbimnNmbG95aRncsTa8
nhdDYUlXVB7fFMlCCXXGIHnRawBDcPuYJuzZNuTqPoOks7x4WVRUpg4etqNwtSoPhyyi8Ghd4XIb
LZY0PvK35gsmCVPl1RApGnDLjJFJKnsdHS2qyyaAujhV2LCU5M1e53egQPZ5gi5WScHViRKJP1+P
Mv6K2Z0zwJ9h5qqAE7IfAtoWwThCiF/44oIocemE4LusqtSU54ihZQcx2MuOrW8rDcZkbDThxhJH
vUx9eUxO31Hlblzy4AqtB0VRi059cxmiHvF4EviCR/qyfFkH78QtFSGAStpIAm1ikdeDIgWsf+/C
kbfEO6381pce1pIHqTrkuQ2ToGjmsHjdekerAvlDrU0ED9/Ga64+0OheP9gvPpp8/ntdyxQKz0Oz
0KEhisJJW7EZsP+CR5mXTvqiDbu6xbe7tlLDfQaOAX/eRt30feD5UlK3ResPJKslhfgyG1rNIxwV
taRPZHDdQSY/xSG21HuC+DCQEy56AvDOMeUzh8FK4ybUv1zjK8eshmIQLxQTrirO6JxL5GaC4gTK
OAfEFa9MMbBiCYt1uCJrku9GjjDJ8LIIwcoc6UyzmZbh1fz/0mdYwFxUP0JNut/AThrZmPBNBPHj
D+xq/xRysH0NnhYexzueRiAgBRwJThdCAcpe1DwWQlYeHKT+rWhn3RN3XLBik6UysTkY++6+iir0
mMl5Zc1M1T806DAd5tRSVDR4s9D04JCAxKsF2KrSUMOqluBbH8AQos4oQS2KV8Ru/QbqmWdt0Fkr
4qcEdCxHyXD0OZdyNAK3qcYxZIN4zGz7+lvsgUqYre0IDumuDU8Zro2xpo+JEEWjddziSgdFdkj0
eVPXn7BoCCEO5v1OWOPmOYWZSKZVlXgWz8u1XRGKbGlcypu1Ksw8Z9kXL2Uq/zlMax2DQEncS/Wv
skphHMbya1sfpLR/17oTFbuaix8Lkx7votI7aC8/oHI6NGXpBSzUegO1OZrAE6CKbpwcHyvKaUlf
mSqD+X8Ox2czRyB63L/0X5U42THJTSoEMu6bf7DDzXfNHV/A5+g5dYwhGKt0C8DWT9hpdhLxujUf
xn+rseM44hxU5rbQ8Gp14Q/HtScGm9rhuCnbInsYs/xK0pMvC1Kll621Z+h2wJceHwagtoBgXvFa
dRha4Qsz5MnDW45o8OmvjqHQnaKatqC8rbs2IAOBOO2Gmb4PLSjTi1+YQKZEBOK++pyGT/m60JW/
mGOl8pY0IybmL29s1Tbx8PJ8SaGW+nMB0Yqu04yL2DU165KlrqxV4YfH74q89RJ5224cTS5wB0yG
+Nk/lduhiKCfKJZAEDmUhgCrJPg4oC0vZkZ6ZC4B4ISmYhtysXXXn1xIcjHE27NDWV2Ri422GsRr
c3XibSdbBsKw8+s1uoYK0E9C02l7j7EagHXNNBtAvVIwKVzLVHZ34k/2m0+9ld02sYF16Aqopez+
QChDL1HRb0ifS1Kqia1AzzIoup+tjj8WHXezknh4P/cxeex3+awyGlarWR5BsDD7QPXc/3x/nob9
yLIJ2IMhyROcuc+aZUcyRNB4BUVWf+zQ6SbSZAXwtpfBg+JKdgMzlGCtECMCHUewysRl8qGJqAEx
4txZ0rWPq3I3anbfD7930E/U/xizsDLYyaz38pkq+xICMRln1E8radvfm0Hnlt6NVD/dNIix/gOA
BkAQrgrSqAby/OLkXIhx4MrNwNKiB9I4j1diOGFvZw0uG2KyqJQxpa2wrF1653A2nLna+MF41k56
2NO7Kr0KIs4rqjBoeCyWUtH+l+a4LhaS1YkHXlKsenxG9CL4yEjdP6HSRE1+wSUnvSPxnEJxOGbj
e68pLOSHVsIEbryOV4I6fdNkoOEZGXIyKr+GkcD1DW6hY1OFUnY+/RwF+4KeBmbTf3moIdYI6sj2
xXUnF1Z7/Bh4CZGgZbE6OeTh+JumW0S4hZd+zJiQB/tWbZmat6LH1iW8eMMP3nqtIzb99N/WUe0l
DjeeEWS5KtGAIBUjBJ/FxQQQTNf28Nfe22/E9l2hELXESRiG3HGYB1KCSYWchz2WCuZU/0JordPu
hBo5gtWG9MuzuubEFpJfwnphQS/B3DSza9M5uddKcszyksVEtq7/hsZlFI6Znl9FFUDK04mKsXo7
2I4oU245t6wGWsaaiBnzpoyBX6hleGmJ6sqvC+sQXbfJiavCepN2EJjC3ulxuttGsHB2W8XAByC3
5zurMaqSCxuE0+atNNNp6s1OTB2v6xrufVBOG6C3prrMQzoe2PWsbxUyCXTCFpgZFoi6ycl+jfo+
VB/w/yoBqflW7zxMp3i2AQSOfABBhIQhM2u0BzxfwAYoo7drGcDz9gA59wdH/9COfPDRc0EbefoG
vUoNmjWS4oDcX2NAcl5aaYJN8XNKLA/uZ95ROXJbwg7UHJyptUctpdHVMMphhtJmoOGjm4jlHTqB
oXdgkpw7UuK6AwiXNXYj2oy1WUsmJXBHTZw/F9UR3egapqdAJHReqV/61BoNb1+Vnenp7rGrQioh
Pv1sI9DorpPLWKLCBJOTr9Lu/IYxDUAOu6XU+Zgtlgh1gETAm8gnUG/2sTpWVFinJMrPnDsPPV7W
5vwzi/3m1kECnOfvZa4xj596Cz/R+OWwDZLbhskICuHYcXY/SkF2nc8zpYshtW1zPQQ88+ouQwdZ
QAuexGAc5LMUUnh619fzji0es2UGNdUEqLsZVTtOc8UJ0mkKqihrxct3PlLMsgjNUpqFbFRc3vh4
MuX6LSbuUH/k4u50qWEmEjkoeQmNJVsV6E4eDnoX7WcEqg5uxGsTEjwng6DhUKmcaNcdKTy8+09h
upcH9KVYrBv5diizVtYfw2XrXHS56DF65oeDTqhCLYTDbtBemYY3OiZJL/MBT2cx5KipHQJ4O9im
VxmZXWxQ6tUUHzUyoUz8IYO57KXrsBIfM7R665LZcZUOKCHBzraZd/KSSmytipjsawNM4ji+GIra
ogvBxXBDtVpn6o06sYsHd1/+mNok3c6IJ4O5xI6nxH1vKf+28FwwPmOdsFxSZVrahbUMVH6JppFx
L/T70DUpFsPUfG84UywE15L+34Ko74vkDuUSWjM05Uwg2JpkFylGepWBCQwSDMi+bHBY4mysLfE7
iDHO6tpFJgt3hmr1y1EgxG7YgY2afsmcwl5jS4VLNX6v+tOZmS451gZebfeOVqsNY3h5ebHvOa98
URItYMiGQxpHpOEXMXK3jhlkPzliJplTHn6/ndG38zpUhV+FMJF6mIQL57rmJ5hqDD8IF4gGFD6B
GotFS2Dupc/GmhAPnvh15i9AEqQd8YAE4uUIwtjU4VHHK0JIL03j2MBA8N2L2LaCfLcE982HISSj
9iBcMrXcuwu0Nu9EgnhMAWuLWJ16ENpGjrEiTuwIwN6SJ1s88caQKTHlacG2gwepwhJhV3ybTIVP
rBmEMvRqru2PMk5qI5jSUwTZNYhsKkShLyp5FoWtGF6Yptu/dJctOMjSkKXRrVDrw3j2SnCkf55E
Oz6cUz2ZT/+uSugdB8aZMHEo20nZ0k7k00AVXhSM9qqMu95J1z5XYI7Wa549Yf7hbi6EdqMrtCg6
qnWjObfAGKtFVh5xrmKEsOeGxnLZtWWrJtQGAPuxp84JeyvNbfsSau5KEdBy0yLhMhLEwSLp6FSI
aF7Pn3TuVbzn4PSwDt1WCsYfg7ntiTfT6+XjOWwfNON12FDISZndtR425byfcqS5B+cnCEtztLj2
FDp2EbjyEOYkvkxtc1X3Mq/3lYtPszmIZf5Qbxtlf9OPVZ+Xd5mx1d9LMEetev0ZuRF0jaQv2T3a
FwEiXhfWlLbyAYQ3rtdOH76Pm+e2t5VwbYmnfuLu547BI/HkT6eZTRdz78zl5PU+nDOz2nmzlk7T
taIxJO95iaK7lwYAh+oJnJy3iAhE5svoFcIGturffC2AFy6HWRxWE4AdDfwKO7HR720nbAk/CPqT
q66BUdKGDnmmsvnqiTv/PfFyG9Z7PdLCihlHV8rSoSsbRIN+NfAfl1xcM/mAFOvUJkZ8t/NtKic/
O38pQV8COfrqN7tZFhTq7y1ORxsqFMZhjT/V44kgAq35N4klChNxWhtTw8lcl6eVlAv9Ev0873+6
tNFoM2RgP7OSbmyG9rS4IzNNRMuwNBQezDZpF/QAIxInlJUe3Xtmla5QI2sFJhb1gIQvr2/ON5xd
jM9wN8LekQmSe7VTUj6NxZnSkEkEZIUxXbEgSS8wihretM6fpSiDuOOdvS9V34wo/T5cUdsCPavI
Dc+/ymB31ZvUcUogS/dhUAA/Z4nX3FK9dWGk5m4xr1tvbm/K2RI99WZoKwXG7WMDzc8wtnwY6bp3
BCl0NlJFlhZwO5SqIkG5ZurEgEOMatzt3AZ8x9eO6HvIurCuXZF32NlJEozIfTttZvG3rNOEDpPL
5Lr43rN94uDb91Sds+p/IJu0tLFeJxc2bD1YzUuCu3T/aT4G/8/juOpJH8Lv8T1amMvNa9Fuay/q
xLq/rwdGuicoKQElYFPYaoOGroSWw4vnTSezQ7wmnPRCsOrZMGPqezAExoj0SXU0fCgIf9s+RwkP
ZBR8h7Mj5leIGcoroC9IqFGhsVK+8zIsciCtH8YacY7v3HTtgbujDiKFKNstik8nbX54XU/9JWZs
wAOlY5aWVPjZ1KCqjnOuE5gaGW2/4mo+ruFriHyF/K+FQV+DadsYhn5ymvFflzRWjpzqIRs/IB2n
iDvimBxkcj7ZRxO8kP+P0/mKZTIyTh2nABM9g9W6qzgZR+6chay50CrKZcdcwZs6iud+J+Vp2Wtj
/SjkJrGNc+R5eyLcxROl5kGKmWl2KWELezWm1UVko8a5+6DcrwzF5R0ufuw4RCMuAqL2w5+KZEMA
LzThm6OtcrQ2y9zHyAO38D8ymHZ1kXAaUqaDZv0eYsFromSjEhHX/jz7rQlGwZSQ4eGPdZ++THqv
jcdiDRxIW39EIq0u4HarVFkjUCJ+hUC55MiCNG8+o34DJxUt4jcRPwMwlLiJ7Ge9dYNQ4sY1QDw1
e+OpiAuKH8yLRDXZCwnRHyRuQbf4uzkzWOtugvCZekXQ8UJ65tjwvf3UhG1IPp86Lw/kkNhg/Ske
d+5jAOpi49G25E/sYl9isWyBK5RviK3dDLyCOJsXlrCyN6VnLyFUxU15SUvGk/WinCmFbdAkFQpH
xdt4hn648cPKJuJ/L+ipX83jyeAtxX9BlcDtzLDx4saYJ0oQGXVnHwSySpn49hwpAxzCKLrWWYW5
EJV6cniaxrosjV9OG4QU4tyU2bRYyWerYE4qNSpuGj6HgftqYSkGruFyMv0r/bSoCSdHY4/8xPwz
iGbaUA6EGBcCxsoVt1BGhGkk+QvlLcEDfDuY3fDCCw7Op4nDkmRVLiODrKyijd04hRK6opf5OEwv
WeZB0oYfOP6e99i/0Iz6+Pt2zd+z+zrAWl2oGWSEfYXHYcXspKeUdwqMvj/U2zMOTgGO90nQwB4Q
zmuBufONkvvt/sljflNMJKyCy6q0PG+KmV4Pv+rsTfgRPAzkD5e+ecOmTfNTGTXbcbX5iI0vYODZ
6BkMOobziBkZlaq5WOQSfQsEaMZM7aV88xCk6eng/myfAl2V62eLfcloyCy/hN0s/WKZJtpslCfs
zwo+7SRAY6QoUAXH4JiIL4OidoEIIMsB1BTJfpvfrYBpx6yAMtOibVN/Fg7plbXnsoQHBSp6cPJc
ZOOELd2lIZpOSuugYkgTCAP5+iPl7+KaypXKb34hxO3i769gUvbuScq5+Ta0kfAqGqBcZ71YkMwN
QJ5rk3aMCOqErBcGLr19Z/6U9VeCDZfraOtXC3lItg7RwBhQhIxaKIxD4q1NAypgz1zWeXt/nCwa
+8HQvOeyiBJa1IfeiicIRUD1pYIOTz8z7C3o1N15BFEEVMKF2MRF8u8cldhWObXc6n3nB90MdTRc
yi1pbD03pdBgxSF12jXhayQhgbBNBkK+g28LiqFG19UoHQ1uMNyiwXj/qLwAqL30Z6GWTxFKi9x/
3LCPx/N6ZFRcTf/M774nXiPniyVdD65MV/2jtXoTD3kQGahxgoO5dmsEOTEOV2OtH0mbWjEG3K/Q
/wurAhe9O5rUlgf8cZpq7qFmYpGOqIbTuLsQzwUR19a9St0IGxMtV+uRikoL/LCyyEfmNNwiy8+E
4enwx9WES2i/4DVjPiNg8UKo2wZvxxibJ6KEJ/hLpCpn9qEpiWj8mB/dkhnM5iMAI08MgqXjkBsT
GN8tI2Q+TAQopjmIL2/PkAdwAvMwJ6ipurNGs4YpNAuDZqGv6KCZPZwSfMF9KBEgeTXWmCPxRekb
OPotcCwPsmHp5CMNpL0mtWp8fObRy5p44D36gxlYo+KV12c1rliwT0US2xqpt/eQjvceoWaJ7k/i
IJCRXj4904HkiGoiCcv+Ze9Mt6BEDF4lQMSr70XaV+k92uKlsMCIEnGOgzUALOm5HdJHPhEnap6j
VZcHgEFOhlj4+4d62dIbp3hzGc2nrAlQv2OMVJdywNPxxxHZZ21uYYYIIRTCI4qrn0y95/TH/vfl
6HDUU5DP9iCJuLsUzaC5p3GNCmmkC5yJuAXPYLXR1VQMbqR/Q2YZFjLG/RMX5OK76fIbHdai7H40
ohuJucuugjlHoumuoGiy8GV2Pi+y4OGaysxSSpzHl8HoI3pkz+9bjdcY5tzkQh5DU5XNPsnYm5Fv
/MNr292HDI/IXLP9snj8LC1/UWDoIH4iWO+fc6TwxIaiy1EEkKV/EPGQ0lJ4heFf//8L+5h8u+1I
CvnFvCLNApLyOQKvvCoGxBJHlAbEQVDk70LInpwIDRgDFnleYetBnSKh6uDCRcbEO395ZRf4/ms0
UGewnAuEpwecK1neNbO1ZRjhI4ADEJ35JGbEVA0ZB9wAflwH6CFXLJq45ojyx4APZCE/uWN49J0s
m+MkBxdr7LcpE1jTjdxznAFzIl1FK2/Knhjg/ocEpjU4SRsH/Ygv8gCutrqRpyUhqvwO1EID2eij
oR5ZiMG4oeHg/Ee9A6XtgxBs2lMt1izHnOmF2zjL6eInM3DSPFFmVuXgEtiRP+F+y4XIh413Z1ya
J16sJQiHS27N18yHNjMgTAwi2Isenr6MRhC7AlyhCrOkrE7rf6YQ0LoyGZqfeecsv5Ymwb5aGaNE
qhEu5pq9IoAddbwyvKG/1ZDtqDxVh5/OEISJDdhheYIt15JnjNpr7wZtj1cj9DPXn4GGqDLHrtM6
CVJYUwj7toQJadLxwIEI4inCLyWVZWhYYQaG7uSvmKJSv1Fc4BhFCe7mOJesLiVWHOa/qyhDAy6k
Kbfb8law7jAUksKFeEu1XR9jHBgztGo2oSzR3cAhfQkN5g6GMduD6r4QI4sLYbM/di5D7wz69qZT
sP5a+MbdxulOM5B1lqqbNGp07OHdJjMy+uoDJazE4Uljvk5wkA1q35SCuyrTknoFnNwxmSLAR5Nv
lr4ujUK4Ni3IUiWS4VYEG1cRE+Q/FuKeNPw+Q4x+TjhC08BDaa3pn3UTiUKi5yO0nkNFf2kHBK8Z
NbdMTluyJegizzKPmRPRTScy51AVdT2TlIzvSMpq6h9giaaUa3CjbMQ1nNLhqPo8VdbtLptzI1ZC
PMKpyGiu4phar5flCPo+PTU97eZ90INawCJUuToXzH3l8vYte0tBmvMZJoUNl0E2NyOPhPMayNi+
bP3KNHwWRzO6cfSEpoKlOZsJ9l18B/tcjDS6xHn0yhbMIE3Q7ZgwxDNthRwkvcKCSIxRodUi+1bx
h7Wr9NHtn68VgJ3j7e+x6KgB7Olt0284R1NBTpOR39PADDl2Xto5SIaeHuWlvRZAMd8JtUs/jCh0
/gh0mR8yj0ByUutI2ow0HTuxorDUEmQ+jCFCkSRy4priH/Kgsjg4wihSOmgAMoKF6wPswqu6QPN0
5cCqJ9jHgndxx5sQ1OX4/f11BbYzVSWP2qBTnpatFrd5cop9pk/nmAT4XUm1VX3n8OS5B7l0kljr
gzEb0AuDJkqfnLSad9NYSYd0SgzWrVqtkAi0TOCMy4mlxDs0KNNg98Yx9Rk9DK11wLjfIuLDvGaJ
8pJYlzthcBXFzHjtIjx5NfeFh++NtggrqPGJ5c3GsRihcLruabEpHx5VMrhkScPkJdOXPYF0WseH
u/KOi1mt55FTvk6OtZ0oAn51SSZjgsbadtSqPUIL8w/gmcKeWjhufVjsk2TMmNiaP7t6vaBqKNCf
aEs8eHPdDl3WyPYM8cdw8cTS4qVuVjHNGcFcsV8GDZnSsd2rZhRZl2z+Aa5YoRJs9fP4zv6tDcN+
HyBdjZyodvA3eZ7saoLHyFQt2OaB5L/3l+Hq4FKxlIupCQEDlYF7RiI7gyt3u42pan77pjOywxXb
niDH02tLCCBXrnLyaJDy5QXXHda22tV82TCS9HO7Mp+xMKraV9h3+gh8cHD98Ayo8d6kTva4s8e4
g6tl3EKKJ49ow52wkTEvLyK3YxjHhCYqA1gXkYUFKaWNLhVjNT3MulADfWobIw/hqWx2kLIG0rmd
JCkSm4FVLiQAbq+ueJ56smDnJ27LRhCoaZf3XR05TiSyTk9OqQ7Y6O0H/2lKVfp1k0GUjLxMFkSf
2vyGSBHdgEZD0c/6SH1Aqe4LR11Cq/yNDjxSL2xBRF1rH1712eMXXLv6Yc+/VhMEjPLvo3Up8uQZ
p8r2HbnA1DHMtRiyAVMGpLHb+HYTPFNISVv34wOkHtUR79wiLSOxQttrjiFcAffMVja7m0oLz5LW
ac/nMQ7fbONKcSa1u+1AjJjrhijHGyOM5cIUCVneVgdE8aYYyekdI16nXauRsHd1yi6x2XupAghM
n9BN+cy47Mw+GJYIdsVH38SrZd/X07WXQKaT38XM8Yz7E/reokZ/AU/07OPFuT5D6PV4mbjiq+yi
87KyZKfxnfv/+c/1Rsn0tYTGlGbza/mYyghE6tzIbHXX2YSZqtbLonv9j/Z+mA/swEv+a83v0DtI
XuAFxU548hnS/LIGcApuPIepmPsMA2In4IiADAjcV4uLW8ZVJ71PkuNxSQvO4AKOhd2KGuS7L4Ai
TuBuR/xMzbNPL9pjHb/VuyyzXJNbrUnx/RYN4/5bNLP50PstYdGbWjR/tdDXif7x4LieL78k9gLT
djv8mPg4xBTFGppjuY072g4LLlz1L6sCOw+KRBQE7jIRMlXD0VBkDM5XXFIfXvl0eegnzUuKEIeW
x5qB4h1Du881s63HsExiHzn/Aet1sMUOW/Y5IhR287cykOmib0FgXQolOCU8e/MZnN7ayZ8QRZZk
d3aFyAL5g3rDQkPpOiaSWJQ7MeMk93AaVXQpffkuG+rc73/lo82uHNh+sSNYlQhyGmrgua0v0Wk1
fPtPPbUEieKtIVdzBas3ifGMncr8Jqv4cIe53QEYWwUAjvvi2LJRYW6n+pNeFz7Yxhgdf+ZawJe2
BUgukxPWSMFNZnGlRP+zcJ8/QEqaR8QmezJlIfWUPoZRolZlAYxEwasqtXK/SG1OLq/egMAURdLd
ncAv9fXEPzB50/dpgubcxkWLi1WHoQ7nDKFHZN3s5NBX+jFjyDAmNy2Q0JWjnNZYFVr5cZT8ao66
/5eocC3O7qsTytK4lJRt0YHu6zSwUlp2eUrzQ9D79Rj1pSxxpzadIgmmuXy+u6f4nLGnQJiAJVeC
JeE0tA0gj3gNolRaWntHdMtxsjJoyO6D4K7z0MnAPaH3kPhQgmvLNIsdpBL8y9wuGbShXDJIel8Q
FNKZw5pI+Q/Xg6uNmEz26r9IaoxBXOmCipHq/Mh1OH8laKFggl7aNrmABMhL57OZrNq6tIrmqAc1
3DLbLCb9EkGorzgf5/hb1WFy8us49mykBFdGjXU0LX12zu5lOvzEA/jaMjIrm09B6jQazNdZZd0N
7oGLtub5idhhBoh1yd0ciRwfXG3p++iBk2twpwcs5n7bFP4Qo4NPyXUr+chi9LOj9IAcXDTt3ich
1R0M9g7XkntF0FvclYbRbBPtWIHq+U92es7X/7cY6M66YQo+G0dwk+wtnB8FSbhO9GLNmiymO1KI
zzBpvtFG7QUfIVZYDNNocoRrgpJ209Fo33CTe2wm27yhbYVAnnlLO06rKOKFWHraCa4lpZhiy+Lf
NbgGNHFhZdWxkpm+4er2yiBBiUo3KG60sbPsU4AmCnQOPaElQc+ZHh1e5sqlTDJauMkf35f/1Hec
B7oo/wn94/oQu3pFvuzEafLKn82F98TBhnu6LPrAZf0JFXiYm6hAJ50Ua4iBc5+NsP/3d1WPZ8Dj
NR2r0NAsRnnaKo9IEGPjSoo4bPrY2haBbi2FRuLBvG+E037EJo3Gvxpim0g79y1Fe/6LaGpcAAAh
D6OIfh6UBqXWzpb4EhdPPIR9C54wJ6Iyh9tMK4Dp6dvMky1cyyskd2mN0CLu3ntd9hmpLUeSEhGU
sKgMO6cin8jcLcuvUygN53/igA5xCk9eJtOcyNjQk9Arc7dwZqoyfA6OLZd0Jf0cl+z8IySFioQw
zGdHzWsbdluyNkAS25aG+Qjx4iBVxyOTe0UZs/gHYrRrkEuudsNcEtfrGknzo6R239nE+noAV67W
8apmj167KySub1faliMWHNv4Z6b5ZGWGbjWrYogyFitOs6A/wF9MakyDm3Zmn4zFEPWRHA+jq9q7
3USOy59raxSjwyDcxJyoMGJzgaQ1WpaUrB2U3od7UKodrKkBHkUHBYXhb+IfdN3B1Wp5yRs3sote
X+Ee+bJe9PPQ94+doIxusYQMI8Z/6jbZSaCx15sScmSWlAsssfwj0mLQv4jDAjxCHbwCY1leq8IU
82PzW3jJ8yi8pKVwjuKps3jdycsaD1y5u3tO8TKuyVBjoKjICamh30khbdazMnbPbqa5dqLvHYDu
LDXGVZcKOm6bH6MTt2FY8K4ziPL/RgzNRB9xIXw3X1FjRWr2LgoxWtS82EmiI8r5BhYCAAcUY7V8
7YeW1F7kzNIpqSs5038UF9zwmgLj22kHFayxAT2M4TkN1s1z0PxnVvkKFfxKHGRNDJ5RtBB7dPVA
dXIC5ikoA92t9zqgj6PN6cPbEa0oE/0fhHOqyzlESyNc5NQBJHafd16PePUQGZXKuSqsBAbL+zQV
nvMGJoslS3oOZt+kkZPOSLGLMPaDPpPC+pYeLLUse5ipNfQKVRUO9OqEN8CrRAu3Q6Ipoa2uwiyA
AmDdo4MLTL2tjAJx2xJnS7A5+V54XwfODMdSOo27VRXXNypslwERkibDywBQvATxcTyQY7kQPQun
UOzZO9rQRhTXCOGS5ac05OdxK6s7sVOSDLYHrEedPS8ZnTjagd6UrIopKXxf6+hDb9H+EPVPHO6W
crVqgq/Bi/D+9gkHpBxN18cmLDKoYANhbASQZgsq7h1n+jwT0kGj94GRjFkyf4l4Fytlvb2MWFQm
gEar5CY1lAkoq6XGPBS39/HJ0I+QS+len26PApwO8p86urK3eUbf1ShGCsukGz1mAEAUf6BF3EVD
Zoz8HCRBmkw8jWFvNKiHkbgWfeZSH0enM3t92tcXvJ+p4u9spnOlU6hKfu0i+4DHKbGJZL4AaWic
B+DL/jthsz4VXehxCfsmyM9AFL60nJKV0MV5oAH1zCyDyHO+0vfsBvO8nxPsXAz8N2F09hBWdmWK
fzKT1b1nXN+AoWEeu7Ac+PSAq48E7cbFLcQWqim/vpjNCWDw5ctLmgvoLSmnuXIv2LQvLvmg276I
3aFegenGooiVCjOvteIwM+1WmouzSlrtPwxMRj3kyWqFCKgPs5C2jhjii3/jGRQT4ciMAyYxAp6d
s0VBP5k7exEs9RzJ975Gi8gV7jH7mXQb6dJ7F+hZwpXsK/4VQkbH/I8NFSbncLNjxh090RgpKtnX
5WLPMbd3ewGw9u+G0JT6V1JlwqcQBnCn7AIDRAAtKJPv4OXJHxZGQThYpbV14FCjAYyRMeJOJC45
ruKxOKc+cIcUiYSNHf3Ie57M7ZaIJtIsj5C/AKkgcN42EOI9KGCqp9J7TVG7ACMw7QM1PUDzhx9U
1lXiQHoyycK9qZD/PNCqACz9ec+GhsS9Luq/xUiM/U9fbuj0+qwgfBDSnstZmJoxLix6K8x/xxHP
aEJloOQRyZUo21qqpLM5Y1WZEP3YWs15UoMy219B4iJIMT6vu03/Sz9hLgnh4XNLMFPcHORjX1ua
f6cj1FGYmlI5saAHJhQFyc/qeSGTSAXGPg2rAyd3COFwiHu+4ap5S3cHsnxVyM3TNQbDkHWDI90U
kyJB0aaMpCF7AuAkHgw86axIGfI5Q0BtcgUDv8DgCP0Egkqdxnx1x0Jcavcw76dApq9OKb3gixwR
vwVETx2k8fCAMjXeMCYjGoI6+0xeq1Kp8/hQITOkoPBgRg9hiV/Y9bBTkzy5ZlBvFOMhTbBvLB5z
KL1WCe/WsQVzbrfyGBFfYbuIKcNeNtS5nk2gpMoGT8PDvLYEYf6Gxvp2l9YmBucA+oAaY1JlPsl5
u6pezlj1d27ntfnUnBEgmeaLL0an/e6DgvICWqDqFJxhRJfUWgBxgo07jsMtkxdDXlxb84nozm/f
j+qVeDakCLFBGZwSm/jwgZPMYilg2VpUHxmCWItGLfe/U2Jj37ACbJmVng06Gg3iDH57+dOg31wp
HF71PTzCW4eX87nzeI0zBRtcMW4dw+URWFx1pkCEDUIK+DgzDdTTLxtahdcmI4Lz0NlA32bhfsho
7QdpdvjIHQQX9T2JPOa6WNn4Y10sQ6as3+z9q8e5gtFljqte4in1RVq07n7ZJDOBMUeglzUK7Vv5
n+tUj3HuEaOQm09Iakf5tpla2RqZYLhrcQaoIAKF2vrL9mBRM4yKTqj9Mi9CPb7gx/ltVh0Xab5d
8GcRf2UJv35jY56JPURBlkJhz0dEveaxd1EJay7Gi3qmqdM4UB/i12uitRQykcBC2Bzrb/TTaGGK
Egno5sj2/UODcIbzs5tS7QlsTZIOGM2pfBOd5TFAAWrn+Mkj877GVw9uuaQuzoGy451Y8L339vsr
XWIaipqnQpgp1bVzPNBdpEa0wtZdyzYEQQlE67zM9PynKYP9NmiXhf5BqMHEHpREcCkFQBDMWxpO
DctheNTjqkgVjIqR53FPG43R8XjzDvSipXsxh9BaSD7unEluQJR3h3nhVAcVU4QQde/xroTj/OF6
f0hSteB+2T4p8ec/79/aq9QpAUC3kQumdzjHh26RMcLTlZz74LkrRxBy41FYOZt96JZuxNjDJn34
xIC/RAyhalvOlHRb+kxdaln8fXfFx/AYsRFvWLBTwjbKTa2/IIO72q0R0TO+lb/WSL4MWO4T8VG2
QVj5B08umK7vifMQE8ny9HKev8ua+2llEhCbzVoMdXvkKZFaGnGhkkS1pwSVA4eikIIiJq9mOJkd
jT8tR4Ekce3h1VibJgCURbQTnxiqGa77c/tGfzKlVO1hX3TgDPm5sarmKNDIZ4iCF9GiN3delNjK
tA9Xlv26ZCuXM+/oUfQQkj3azGcsSrVXq0LJ/kGJXI8wc8CZkcYRzF6XPhDncDMEGeK1ZtEp2oKH
cwyMB+ETWBH0yn0uAKwRd8hz0qc42VLv68n2ev38UHVdBF0EBxpLwwnuFBFbLNwACGaeJ8QvkPIn
AoOVwYpDW7uewP5KOMLh34Mm/WoCHO+mibNQlsTkuWSmmPfNhmIQKXZES6do9CgqJa08y7RHomGK
KNouLKdUnEE8J4PYXBzoiiKLg220KuxsUibJf6nRuNVMsvy/vEQAjNIl/opuJbBS0fp4MG1mxDB6
GjKSfUTR1N51p5fdV4Vs1MD16DYklHXxniLB6u5kmfr8ab+bSEpdeoMvjiKe5bXIRAKfkv0ouApk
WJjgvAYI+sHKS8jeFxqe82Hnd7NiFpzdJb0HYL+KlxBja3E48so6V4Nbdy6lWACODz48e604KpmU
/DyZ2c8jj28gmFlH1Z1VCBTcHINciecIglk+W0wbfyLr07k5NLpPdOBn2G+zF00gxiz7y15iai4p
mtsF+XqGsOD3DeCE0xQdUP7hgq+eGjH0470chhe4Yrv6/PtgwlpaA06wmkBY30QkOOrYYau5/Uo8
CIL8V48dJ8p0PAQaIVHCnmJN7LuNOohE7PbC+24eRJPoJRYe4/9Z5uoCdpzuHL80fLibhfKxj9xQ
FYEi3LqtfCc+tgEQrNkGnnze2Z+PEMOFnUWjDtKApm+oU1AgjJvV20Am10CJT9o5pWyDcZ+HiNZL
+DoDoiv0eCzQksMcmf1IZQQGZT21mLOr4EF0qo1g1E2PqOBbsezRnO6tqfavtw2UIsTCqrHiOIEg
xpo9abe2tDtQPJgPgVhyqrGdL7HVm+F2F6JppCu2k0UlyRYLk5GsuIIqOv+hgvXDRumcLmqEmJfY
WROTwyMasPGdTTrEZ5J0zMnZHEZpe2wcGD2i0GZzgf9Xc33QuMSteICPuu2+o6Xei1CUk2EIjLzr
29pKfshIoknj9Ms9U+MjUTYrSDcxLuaFBQUvQiXE33sxuUz9RWchuFW2i4lKSNBD8uO04tg2Ct+m
JqGG2/mwJmwL4KUnEhNY7rXeCO8oncQOyDVJ1JfCRcu9wKpuvIsa53RalOmWU49D0sw0p2pzXwRh
JtCloWXAqBEZ7c1ey/ZX7kl2CJ5k6C9JSIKXe9RVBjtDoGicGqM4WesM1nMuZB7OrphOSuKU52lo
tYncUdKfCSIpOn4bLhbjigiYSWrLQhFCfymT8kG2PEIQLPzyTRiSQlOUMosksarX8m4dcGk0jUPF
9ZnZUIHivGiVwuskg393KsxwcFHLoxbsNVQNx0XrDx5xaREw5Db4mPe8f9aHLTD1b5wLHJH3dBtJ
cm6lwQ8EJO5XRHqWV0Wel5Gj812kmiZ/wBK8kPQhsVh82RQwGmKd2th/JlKQx29duwl5bNia3Odi
StdF6TtRfjPJV+D92u61UB9AjaQ8EtnGsriml1suPExv7GDWJ1GqMucf09QApmzq0F80FAFp7zt7
1sKBFspQs7f6nOfJRS7GSKU/J6yd+xL/CjKqde6OnzzL5Za6A9Vtvipr1oOfcK2JlCbWUblKVr9P
SEz6k9wyU/F+Bu/RKBjzDKYcsn7LTvpYWe6Dnnck6TkKWZJ2H376Oqc5gZ4EixpnFRzVbl8Px//k
gqPPiBiIRumOjXUmjsj5k1ehcUIUmlIWj5fDLnQS2L1ndr++fYvOoxjjNenM3zOhONKA7//IQ1ld
Ld24oO/1Mofz/LZZiPfyu/076tZwWKhrl19PMkmQTsDB4a0Gd8MtgDYftFqRpNu4Y5KqigCgQ8nV
XyLNibXZtFn6hqhKJYcdO8jz+STEJg9O7j1Y1Q6OVabRQhRZfMRqHym4Wmu2lQuDjBHenA51zCZy
aD/z3tXy/22LSSySXM5oSuH7nydxsUcsU3cQrILcwLxIJTg5vTBx2cBY8Znta0dymtfGepTPj5ks
QezNIKTLT+rSU2R7mpMUD44lX5PrLXFNCdsgBQGTmPhrx7O60yLwZAENE4/lUnfbBass701l4YuO
5GDyV1SiLmIp2Ad2cMze66ZZcLCzgMCO6rAJBcRbSQSEcM2ulvCh0PtgtdGw1LzX1PK50zG3Fjd2
M/a74qFXnWCApZARFaJNyRyzAEiGf0ayZcN89j2Uii6wKxKWV3TVhQ2Yk+gDKaCtdIPVOfmV7alV
51zXT00I2Z/tEjxZuWLyM9rccsT64k681R7xYf6/bqq4TNNdhVRvDaENN1eFeNWCzv64k4GBlON2
hAGssFuAL0iONya6NkvyHj6mXGnD7WmKPtnu0GVHa3xm2GiZW7A2jRTGsttCnz7CZKGwYZc9pAvt
2re0OHz7lW+0L2VvAAR9ub2S0eb5Se1paDjQfZnGD/4OUqZC4KRY0+OhbJNed/JBezZE7eC4zFX/
E5QuIjP2iOdCf9aVCUUMp08gZGgQi/zKOhOmPKLmIAj0haO9XidnURw50D41MInpIijsqCJJEpsQ
LWFzy+uBrKklR6Q5/JD3vhPwD9DXEG7HPzm6qLU86eiuN0O5kt+HPqwcpvrWIzWY0u1a2ZudI7Ih
o6BKaqsInEh3ehH6wrPRAeGOiK1sl53lhTPIYt8jlmadlC2kzC3IElVZnQXkesVlutmei2QZ+qSW
gVcHimkxiPhpWbKTMHOygg6vyXkGzkuI+3/KcBg6HAeN4ePbaxqzhFNBmXAUZnUSTm5IYbHBpW6Y
PKqH8MsZhpPd44mXUX/HHsBvqpypGP0uDqrZNMqZVng7rnWLYQC4eypj2LTk8iYms9+Azjn2YFCn
SqS+6P57V1sYY/KRW0QpdCd6mes514ee7QdEa16QyXGJE4PAkDhmqZ4k4sHGHZEWazCtyo5gQti0
4Ku++UnWeoFWv+C1OAgQEMJVkaNZNF1CU60IPaudf5g/UbPnPeIBDYU0bQEyl/Zw/U1EI7PCMu/K
Y/obLM2cSir9wHhfC84U6tMQuCntYlhXusmbeLLsgpj/lTMAbmKlJN0Rdfq5o2JqoG6klv54V8cw
6qL2ochs2n5SeYehYcGizrCX2pDCJWKh+yfCmwioSjZ7cKMW9CoECOuvelJNKGl0W3XvBAknQoqg
FAkdc9OMe7LhivF+cCVo99vuvAtUQBED1qrR00FOywcYWvUu0f3+qPkKYcMqa0o5bwyFLkZB3GJL
AGRAe0xFF3ZJKv+MdUZftcW6oPokoDSmzl951Ebgs+DTYRXxT4rLteEsfk3mylaoiMzaloQv/2Q1
OWFgmuWw2XHhz6ahaRPamxZ5+vXNjYNsO6gasFuOBTn3KQQiqkPf2Wy6StjpUz3Ctr1OLOluIHro
8i+8naokcJRvUw37H1JbbWStHECOdzbkID2wp6QspdnIoG0MwQosPvEbKZIZfM0qhPQE8BFqydGK
1Flyq3fizjpYC7dsaJyQwvtui1ThuPkIkHK9kRaN+C/vmteEe69dIWDn7rIIczAb3PyU2VebMm1h
Xcp7qJpIGULH5sZ2HNls/Z/mhm/rEleOleZSPSXK1nZm7qNyP5rg8BZT+cLy9/x9Wjkgrfi/4uaV
i9heTTrIlh8BS+G9MYDDM19V+58Sz+2TPP6x/3xuGDALh/MTkwpJ/rNi9gmr8Zefyczpf4aS3I0K
z0x1t1VugSSAYSSudKGEuQIhxMuYvX/RFURzJE0oO4J3Pnn4q20MXaxzNXjsIrxGwTWtDPM4ZwWB
MiOg7Y//1CtuBHIu4sXZWMuVh8pHBk4ORJ9OeslTnla0eQk1eNL9rXLfsSDFZxZZ5/xwDDqwsB/c
l1e7m6ukpfnhhpbQo3sFkwzJIxlkAOQgUTcOrQ2g4EKd+jynhJMFtTiPckzzMp08CJ5xm3c0idIT
ZT47sMXONvCGEYjTOQ7EaLmP9htFrR0kbXIdVgQu1TxQhkjSNV78ysQ7I/piVauBqAtICn1GZ/6r
DE2NUkSryTknPwhbVdegQZT3tb2d+CuM7/JBZuhg8tWMdC24M3sae2xqhQ84Xh/R1pqMESpneRMS
QQ8wV2EvgAVyVIQs5Nlu/9YjX9p0OJBLCoGbIk3nw3RxxaLhOwXKV8c6On+hOEqF8UnyD+G3tluX
hWs+FNrJXI1qvf5XhD2jKEwkbsFB4JzoukQtWChzVUSjXuinbLU5M+K2xgZpTsbZ0PTXbef2twCA
Ia2EVe6mOJtNLa/pP0oO339MNqerEbluQTlKq7gorHaWsXAaHL472mEIzA0KSQIj9troMPxax+N4
56M/XTfQmFdp+9OcG63IRD7o6Ra27+LhK0hmdZTAB0s5lLHpiYQnrTeGL+fpAoHvnK7BiRFsRw9F
nKupLR5reih/EnRZPAwCjhlaBSD7AwiGsvxOsZvWtDLiIuPMbm3GqIKPHgMW8EtkGCZwCCHDWWQq
huZ3YrKKLeyWQZ5yc9qmOte1UMerbYv5dnNJRgi5jTp8+DcWaciu5gVtfKKlG9cUlQS1CyRBxtAR
Yshcm23CzDc7/fejrxF6UCfuNXjNsaakSIYpVDH0PG5gzWdmZDdj5KMjAsT4c3wrLK2TQBe2pVP3
x4pE6SeJ1DbOQQAZf8S+TzMqNc0l0xK8SdO4G60JFM49sHOoPpoce54J5bZZgjme+wyxtBZaG36S
j0p5c6AWI8qUc9kA/0fjXjTEJEqEiwRxIGfxnK1S4N5k99/rj8VL0d3FUN8qThy3brbdp4cJa+4+
3WyKN9J8y1aYKiT/4ShFdUyueitorBK7jRUU/6QAmo6QOefyLzax44BPguTdCQ8aN48kDOQewvNT
adPoBztMUUsvz1yHuWp5/tuVMkV0X8EaZl7f+3F0Y1sUS95i7uo2CBtJ6lSGkT1hSSR13zVP31F2
h92Z1tRtaN+Ur4R/n9GrUOVcymfcpPngFEEbMJP2vJbMq8IvGUbbIJTjiSJlWjXt/R7XIh0BASKE
OzYkLhPF7moXmDj3fHchlRmXPjBB3gv5zfRw25nni2a+jbp8cZYw95vmh7131lhHKbMq+un66z85
o9DlGrFUE5sSuQubG97jrTB2fSzA8lwE5JSaBiYTU3HHnZi7lmtEpzgti5uOtntz7ydesUo2VnJf
65WBwCurwDFQrc4Ggfk2rQV8quYnJh+6lHZRSe9+U9SWfTOU1dGf8hDwEFUYWkQfiZxeyrHcC7nC
kuzgUFEOLhaqgTQndN1i3MD1poMAE3gGzoAwZWyHbrcfUj87YSslW/YgPK/x/g2KAlHm/RGeflYp
AU5FymeItVjsNZ8CP6F3N97qj+LQ0E1SqGEBCLJltr6YSL4cqodDDDFLdsUjyZJe5+Cwotz1dqYr
OuGgXIFnp6QtZvOIK4aXCt6u77BWlng8Cj2BHCDCwuo4Dic5YmLIL2EnoYzQvO8GNPfupZ2EQMgB
VDxYC3KfisYjWWXmB7502lM4x6NutWqrtHWPdvQ7rqhnA951LtnHgfAr2iB1wQ37Cf4ug3ivEEhG
mELmDUB4k+mQZXw5VV3Wnm6C95c9mAx7UVltYr7vFkuzGS+VvQtIwP30PgH7/5BAh9Dzlk81Gwys
GIBfswRv0eUfSLfmca7A0E+knmGMSvMzHE81H4sUL1f2TcW385s/tloKnF4EKQ1oJghxj+H9HnuO
18TSMRHEo/njFmZmR4jVi4f6Y+ofjSaW1G5TLYjSf7izS//MKl0Tj6YYjPjEq2uroPHIGSzcJSMc
6AUI3JiEsABTf6eC2yUhV5FH0ZOIL+9NxRFDJOtn1Z+YK7r+tOkNg7exOvCk2oU/V/HExYePSa/1
YhME17eXuKoai+Xrf1vXUCstPBbKeW2Snvhw+PzlwZ+nM3JwOHom0SNlg2YAI330WVkduGHa1BJj
EcIIzeWrRXfDhXmC+eZU0ZvY9eS+GkTtmktqggtuOfbEd8fWQcQVJKxEEWqfkINjxZ7RXX2pQ6kB
+sfQFDPpGdr5Ld0MNHWgtKX9r13FwNz3cLLlF/MHptPW3ZvKpNU6SNETaM0OLhzgQQCS5BeyysZS
tlrg7Yu4ESWyur2uwquMMhzRAF2lZ5wOhs7/cALnPD2rhjs3Hfvbu7XhoNkWnmLa4pqhhB3/W3QF
55pWQm1Zv4bWibYcuSVZwJecdL4FTIwBHnOjUA/bmzYUUcW7W9ko8aCiVujXh3utULhkLFrkbnRU
ovcalz31PPIvFrZFUh2k07ODoMYo1874AiF36l4YUtSaiOLrdcotlWjR5+y9AvgASCqux1j62wSH
6BcOUtOyOWFjVF2S2hnC2Cp7yKGdVjVHrk3WhfBzhaTSo7TxxA5jk1DqfhJLlspSKf5G5hitqjJ+
oJ3EwIflKPeOM8xOKGVrQ+4uQ4mUIcd2htzZjIYauzvKfG5TYsYVAC4U1AwOUBdapF6oEDhuESrd
mXIrJ+oq6sQYr6bY4P+vGMvoOCDWvgbhFYouLo5zzb+nYeE0Nfwed+6RXlDib7hoImue+BKCKFnD
S+rkRGCfWJQTbYdvaa/HZZ+p5niu5lBiBpLHsmPhLrPEDTns4hfAfd2yL1KJDyRNSkkYY8f2x2IE
IwmzYK6ctte8H5eJKiBdYwIU2h8xQoKiVF0iUWhagqz8rbZPEL9d7QDswk0Wm+7JuJDDFXx2N1As
f9ZicZ0P0cW7DrMMi5psB4mgfiCLl+Tx9dCncf4sf7J4uKS99AoIlAKodupxpGLEmvubvC68fPu4
DSVgUitpIgsx3hVFDjDIAwEH5OtUOAdeGSBGT+ZDwxeSW7FCuPAQY4q0s+OjhNFaLWQa98UnqUy/
IiJklJYQ0S02oE1sl90qLH+w/vV3UKHGUI0AFeyJW/qtYt9tSO0MxLMOddEjVhb5LJB3wWYHF5hE
5yzTcmGim+6zg6QaDHdNitLuLA/VSNKrkZB2y/wYzsLTkbgQxGdanRgnovdLlO2aoTGXOj7usPZo
DDLJZpWHbHaG2r5HQizB2nvfZaacrZD1JfnMi9v3t3mMno776twkQEjCg/XzZMFOehP9BqwdGRdp
UVkwodQA6gEIBrKu37ScuNaBdai+NQi+XmNAklMyARoiE83XuDR1UKJJxpy1m7bXnCCLOdaiaWpQ
CYO70iM9ArKi3q9rZKgt7n4Wxu2MyGVjGuOo2J2yb3LgS1w4AitkF3v+9lY5UwADV8lYo9aimMEg
kiG2hOEH6heQIPo3ECwxcCDUpZsyKq2y2HGN9z2INzR2J0AW9XaDvO5M+D0B93iIZjLvUO63/9au
Wj9N3GsLdSpDB8Op/iU4JLD5tYvraLPxjh2O1rO2g7gqFy9OYgNeMBYEhZgWl6o9C2DedqfCRob/
5knCqINzlyctzM2p0hIa2shHUD6Cq3z2LOUdn9UzeOG7l7WaHkp5e/eH50bq2osbv2xfVw2+f7zH
F2mwdNdyEnIYLMAjMhsVOqP1P8V6/BlhQfgkqBgEftpnmTp7/ai3R8RYgaFq0bjZTO4i9SMvEjyM
DFBCu8KAIfhPADO3TSzu9gQ40YvqxxNqcy9wal1jhP/E5FEDe2VSHMYdGrMDs2rXbKPqmmNjeHb3
CgZktgBMpKwlTTcQzh6m4SQ4Xd0E11OmKhnldxCqcBN5fsQpGreFCanC6n7E0jFsz+fGAcaSCHz0
9gwjxHI79Npygeo0CaMcthMxT0LZjobUw300PN0MwBdAwa7bhuaSwuK4W7ygzzWYx5lroed7sPFx
4qv1El7mLdsoypR9fi+6W8haj+mwLNNYoMu6828wLwG4WnygfqDIR2U/IMB/0ioqEUz+WassOjux
wN1mASu8UdndQ6NJz3jlXcdVw67Uk/CL8cH2bezC4EVwz4/yDByhPNmo1ScdGu5tvzOlxtun2ZUB
Q1Lpu6tBO+tbpNcxRFDojWfSdJisyx2MgVJ5Q+jzy15IDG2BDaHBCjJop1/QGNj1UVdMS1icpHDK
0SWzH8ElwYVPNXGH9vgobqjscqeJ1uGwJQd7p3akyVKlHAGmVBW3iUKFNzJW/nrcJJ6LUccxlmyG
arwnmSY4M+hupNgNCHLqUpPdMvH5kL+dLS4uP0hd7KxGhyEOuLYFYuR0bMDicSt5ObESio6bm5SX
snL6X3ClgqEn5vspSakIaSDbpBRTeVcbW5gZ9al2vTS6MWd33hmF+kV6QE589ry6ZH26xiORFXj7
z3Nxuqi2HgE8HQWncRXRWdl4FKhIpN/aThmAxq/1Oc1mJXdNJORnTKw9YpiKxq+JBLD5doLECUTu
UMWKXACHOz8k+gQhLD8eMNwqURERGvSKPxALuR1iY3/sPtl2Lv4tyxtXZReDb9W1fKWQDxrpQ6c6
OD0R1ICr2T+F+rbwLcQAzyvq+y5l70DLugERj6M5cnJdZE2j7/8VJXF+CKbAhO4hSlrWQkbsuT5w
RVl/anbIArJx0u6NugzDz8d1V6s61HNrWTZ1o9GtgmVHmrB+CFfCiponerVGYRwP2N6BhUzrjBy5
XzpUESz+vuAP1+dCkBrwBGvvw3uMWvm5qmp6+BTAGkw9AXTpcySznA3pC3h5ptL7m3jb/r+dA88Z
GD6rGywwKb7HFR2ob3RisiHg/X9iz6c9O9MhHmZzULenX9HkGyX3j2+Lx1KPvgaN5qLWBS9cuw6j
eqo/pYPjsLbTdS0f+2MWezkoDCXUkhpVtZGgPbXmu215KEyW0e9EmJ21MVGAQZWmhAPN7IjD5wn0
C+Y0liryZMNxf0y/HZcsxp8vpapEd4JCXa2NPzNPnr9K7s7NDyI76OIEMB0Z9vUSw+lt/XfUD2eF
XtUBgphU4LyB0hAJneOqCoeXrUOGFKqPqyo/oWGRLs3KvpycEpfqux5ZZCnAYiXfoJCvNBNRUgHH
kQX4o9p8T73IKWn2TkhR/9+WzASvcD+VQzWugEbBXbebyqVNSKskHeLkd4tWfOMhTFFr42CCp+YY
613GXrciNB5fJoDolZzgRU7jqmKGjLW7J7uIN+urry5ErSiaJrVmHjEyzZppMVQAhu3f339bzdEj
MVjpynYy8RUA24/dz9VegfTzzLhodAuZt7wHyGCGeAmy1eWLJmFJrZsCTPEuulJkLahQtqj0u9ja
Qk1M04DIvdieQgX9g7qv6yacomOugyRK+mPRxP+wapJIGRcr6N4H6V96+x6PIuPuT0d4G9al/OzH
9B8+oLVr+UJQT2hZXJ99rm7P0xhueqdc0SDmNA1Gq0S+RmyIfsgHl+aDZ+EX/BrhN4Eg3ghD2OV4
/W3X9IwNUxp3qhFQAKO8UmFtMhd6kXttvRI5k8m9spM/iaXHnackOM+T0DfsqfRPD95VbcIhAtRd
lnOUhrgzyHT0oWrDa9FcPq5GtpzvaX8MRALAHjOofOuJBK/OtF0wbveQH0Ot+M+7p3FQ5+2xzKFv
EH31ih8kjhjny9+b00aTBsn9sq4dcDmhvvcif5GOMGW7Bhef6hCXjauLQYaD7eIe+mTFaD6SccTR
/qcc/Tbfi3iV369ohm1b2Xzqp9Noqj0F5cfan9ugTSMOB36jEuKcLM3+2IXWfEC0ipc68r5DYsMI
THqzXuuCl6KsKKuamYpaiyxn3pr3dzVnyHBdOkGfjhbe3igbygD7sNYc/Kdd+K/EQp9HpVRMPpA5
crZblj7Tr08GFNGLZZgyzBa94Gqj2FZUp7r3iiOLB2eaQbfdt3k09GlrOdhDq/vNZErkGMadKQTg
StPFOyffiyeGMn9PKjztk3UBfY+Jeb+0TEJ3/lUyuLhYbzw4EpWpg5UyZzLRh3VQmbEAqajCLivd
n5keAPBRce1M1ONPzi/qPnaFPC2C0IDTgTTULrJuYk+LxlLs09AiXAp6lhA4I1puXMSlBrO6/NJl
YxnfVlK8GuzwLKMfm9CfY3Z3UT9g4jI72eM7v/VYxasuFByRWCJYiZ8s2dSqTcxoxt1syqIAQBkK
qhopeiGD/9bH3aDgwUaACaUa7A5WJu+7qK5eEJwKLLATn5i5ORrUPUlynTAmU4Jz1utbfqty96Kg
6ua9AgwQQcuCDf/7ypngXD6FDV3x1v+chaugFy2Id7LdA+v+Gy3rRXHSDhyV/1dby3XgSfSADH/V
zfUvZy9GONsngy4fju1giDuKqprUsK3czLWXzkCruLvQqX58hGXzH2iQKp3t0RSnKWCP30eVd/hV
c+QcAz08m20QgnezCQRHEoWPxVP8ZEO9AIlDmkojEfneMpO/nbaNnsPMRVmTzuc2xrHabKBY6P72
vdvCIWfo3YGdXmTj2HYDGNopddGeGWSeFzy/Q/vpr5HjeCwB4BMBcFjWKZ5BVKZGPlas73Rj9gt+
reiNMvBRSCSsxvL+4xPRd9u+115wY/iGVH4LxWC6GCkK0TmtFgLa1KlKCl2wbiBsjpZi5B0UMr7U
L6VJf92yAMdCODUQ14ayGrVosgWV+XHpsZEVFa1aU+w1AHocPmVfCfEKEBLU4pORFdqu5NSurgna
xclyXlaJzowyu5NZJ1tVX9NvyKASoIaCZ0NNNz4NEWczGKmu6kZK8SSuGiRPd53jyCI+lWC9Q6Jq
9ol13U4U4313D9YckB59fNxG71M6OzA8VAGpjJJJ4+CWKEFHtZr6uUlSn+TcZIBkMB+xP2RQK9TB
/999oY8X60Yn4aYnIsPYUKb3X28QgR3A51aEo6KQWs0MlIydQJjV5f+8aGQgwKF/Hd7V1mq95bD7
feRW/TybCR+hJqLE2SbYQD7uCKTQl6EXaBfBoe78+ynitbiyEnGImEiRS522KALbqbfq1hhBJ7WU
+E+fhtKDKY47ICoj1QmkvBs/mm7YyyWQn5+47Os+X74W4EMTy9jcfoU8pYngikpwdO0Uo3R7EBux
cEZogK9E+bDffIKqZl1ZdfhoZAbzgx7mFYlSQbIHbIAbqhDsAdzuV9sk5pmNJSgQLEH4zIWTX9d7
tbtwWOqvKd6cOMKldu/PejfsaaK1wAYc0mL0ACIhiQhqyUfh4AK51y4HiSY036AekWTxEfxXC56/
g8xW4nQ6Rsebu1FjzxXZB84BxKJu3lGi695efWdiQtxOUJOFuYdF+nkemmuuFFCtW6vReiWCmBH+
6GE9QIfdxHPcTpZGmSlhplNJA1PhLeJBoNuQNhobqnAcjlHRzRgbyT+Md94SP21YW61IMiFhBsTm
IbNldRtxGyeGFmqI5F9ymfBf1iW5Ori8hMuEc1FU6KkKZTLb3kJQ579kLfG2YEIg+xVGFurzdZ54
hwsamGZEIYpoCb5E8bElzRnoJhTLJSNeZRRUTY6kodIeem9JoV9OAtyPUQ6rYIErJ1UiHxuzMbQq
MEAZEo9MhrqrGnOVb3WDMf1UCjItAE5CFoQt0F44ngxdgEmTlo9W8fdf8VUgFHv9OWF1DsOQq9SY
t4zbZizWoSuIsYKa31gJgVWjhAB++jWoFE9kWPK5J1gB+x1whko4AYZk4AFnwwteE+sE6ECs5aj1
pG0llXk1OAV03XypHz/EclTIzCuT7g970knFS2D1ZfE2p7IfcY8vMpxoC1n7x2w9KVOgaeA7ODr5
VoqQfBPX0NDluwPBq4RJZkzdg+u/K8s0bvBz1YnOFvQzOS5fnm2CrmkYtKrWHTV3/lQwZ3cWvW8A
hPIvBwM4e6eXiViRNQYleCrPo6Y3JX2VoDGvmbg38cgEVQQuHwG4KwTgeIJp/LdeOyiuTZTU5lOu
Iu4D6IkacwjHqZdNR295Os18/BBbB2XyHyleTHI1da6V6mBJ+noohmtUeJ5PbTogVW+i0LbDzSUC
8HaweGdEv4uKzZiwfi3vc4tthguRjkrhaot+vBbYXO9XIhmjV5Q5BW+OlxitNeWKjL2MxVM4kKWN
5vk4pC+iq3Gq+zokGvISA18l4vnC2HeTLCp1yv8x/iOVDN/eLC1pnRF3MutPrdzFwhGy4qEoFxe/
PEh/BwzxKHXAjmzN++bSDtbptN9OoqqU5tBYB/KC1KDtV1tjJ1jMKVxh2997vWRuLUIWt4TkT7Q0
S5rrUO5H9fGzBeOGwtn9zup9HW7j6PglcXwwHKwWLHTSjfGm11quXygAiIjtGTOKTjVJJ9PhxGnA
oN1h0ucc4E8SHAwKBejb+qKGD5PfTlA+haDqsJu1V/SoJE7ir6P2cPvgfJo1bd6vRSTxhTa5E/B6
UtKzTEbvGT/PwD3kxHcci7T1qJfyQNFJ+SGoRt4m/6xlqy8I2zHKVVdOo++8ixS3Ab7uWi/31Q9U
0UR8/YYBvhCLf0mhIzYm7SSgeP+Z/LAwgsZ+C1dmjE46qQFteBK/72BK6/meDSdh2RK903KnQCHX
BplfNLFBbyDpOS2CTxhHeYAQRPTFnrUQALzXot/5N46cfVv3lucaSvHx9TmGtu2Om8VBWIt3GOyp
9+kZ7wCF4dc50s11iTNoyMDpKwCWmlXOChzbu/B47fjEHoLQnLkXghvCsgcvK0JUodt8V153ptnk
31EtKF4yRAy5qggniF7zpm7LWrbSOzQ3a8oOHMsH3BL73Gc2ODQmsj1AO1J0mjhy6gI1u/e9S7cb
pKjv/R1F2gx7mpvQDb0ZW7xnm9Lu3Kf6QOeVNtC+FExsGgs9CPID1jRGO2jjyXc3seTHIWhyrFwv
ASW+Wx9z+E5CVVDJOUefr7Bno0P4hyd2LC/KiJmDPOA1vZcGaRmW3hD9BSd2/zJ8TeXFAtgg43un
CaEig6Tz8EO2gOvQlVgVKAYjeS0DbqQc8du+kV/LtwMqckywoIO9k5MYDBZejUFno1CyMiEnqZJ6
GiRBs7aXy3/CUFWgYaJavivAupGHFof573ALh4EYA8loamDjuKnNi6BiUiUsy14fn2F1FJZcxnRX
inVTgTBGlvltZctmVSKTBaGdD95aPQ4lD0QQlUEvPGT+UQZ/rWt71PUXQ9YXrYJRcIsPb4uRhFc7
S40QU6ed+PfjOgBio4nTLaLblaBPakgtwVbTOxo0x5iMeH8tYruOm5F65TCBPBMcmVtAvJi4rRae
XKQnAJf+vvp/xfaeJ3ActuioelmNOKBWOpAPC4opf+Te6Lw/Sr3BpDWJrUoZYYomtqmCDxEYxsSU
YFCUN0c/DuZ+2c3TZ58omZtNcmWDzik2i5rTCwEs3p1aRlw2wiYDk1Z2wedT6o9oTXJQ7x6Y7jpD
muPm0/rKD8cZt6v0+55E5fXCWbpFMFRKBdYWVIKyssL7uz9kKpH7G5gyJ86k6TTDmFwjT4WL/w6Q
8lfTHyqojtMPRyYAEWTEL5dltaCMSatVOa3FsNCGnD/tXag+/+r5pQqiCYHdutPKB8jUiHy6phSR
qvJCEpp2PTG3EwxLtaFlQoKSrB9UNGk2ovT/0H+YHVmBgBjfOL2N4QtCnzzUH/4ArnaAwrtpWQd8
3ludTpunGEVEqlM/vZ60s27t5KULbJa27ZCwzk0NGWCwHLbhasH70DogBqbPtn0CIHJ5LjIzvvUG
FWQS3UQVYzZ9GhJQ1kuzqmZlglM9YN7Fzok7LAe6Vo4PdlPvxIAbN0dR/ZdulzlRXL481+O3+2vr
SdHR2tG1trUn8cJEF3AKpsfqb84c+Z9SwgFuVhc3N/KDhKshJBXWyFz+lyQU7BFENBemUmL84A+2
Q87UX0eobotxTsEpfexEc8NPOtQ8GF213PfLNWJ6niBV7WuA2pHWiOB8N2kqE4LhXxLlDQ7BRnEj
qlY92p+MJYRG1mTH0OdtyS5aYS7NSB5GphIhlaJ9CDbUeA18gFTXNhaDOOIFF9+Blrx2ilcf3no+
ktgUYk8BxW22tIQ3j7UQAhTIa2SdJqwxIHXDUfHorV86vNv/GLAQh9IIs2tOwVc9ILUpGGZwjqpQ
J0KHJ0wY7xsOxKy4As0x93wkYkyM7f0OgGQBhhP08e1EC8TGH7r+Oii4xoPHAMhi2odtlSi0v4/M
DDTtJxKUjZHljQ6ta+qpU6UCqXVvLrvidpjvx8hDpR6UjESvYh/Z7FlPumgKrwBr/+hwSd05wUjC
fvclGZScUreCKVqCFdoR5MPJDIocPDb56BX9iHofd6szJfuP3qJZQohmwZkaB2Qwhhwf1/kNFwBZ
eOojxuYELZUHG3FbQH9rD0ERYLk5pl55pliO5OP5uDM8iygAZAwxhnbABRe+Uh10XyULBk9qcxOA
tZm6DfGlDKYp78hC/xHw50nPTe9qU0JL2DUCF1ocjPo6HfZPAAXg8jYGqzHPZ0QRAK6SauDgkNn7
9Rn98Bvi0jTKtsgKpvfaXGucD8lOfSjGfHLhY8PvyFWwiwoKRhFPHXhSl9VF9NX1CKMW0ksLzoKd
VvuDyHXDy7JNZZ2DoIL8hJoex35uaN71pvfE/TWDawfkGRPWvp+enEjRyCGJhOhbnbYXUFQjLV10
t6a7Fg2WQE+8gx+i+pvio6BIPdiZoUGzqURv+e5o6Y3BnBnZiuyREEnCXleiuL0GYdl3THn88CiZ
LxdFcceUs5BhYvBh4huaPhXvoOb7p3+Dwl7Q1Qc6PTIis20iVHDHX46XfOaqsTGFIA9/bIOEWDbr
eAUxB7tLFeM32HZSNqVydIq1Du8dPJYamBSk5II4u/wXV8xHawUEzwojJXwK5pxslcEp5sRGgxUB
4TlmpO4eORDthM2YOiN0GrPuSfTcJwFQP9kjXCBDkSGC2p8Q2a+6gFP1/G32Zh1Bc2loIEgmEVhG
nCW0OHo5EVarU/r93+Xhvvgu/uRjr927AIPXK4+J8kOEuY7zA8KoaHg3+G5CLcjO5a4K9R4ezW+m
UI7KQEOM8uRd3U9U4DLUryYAZ1clHvASE9UCG5rAp8P/RPj05/cOHUKUXbOkuzrCxFzA2LeS1JBq
Fx9hZ6/54F/thp3SPgVu1ye7trVrvLn1UMo3ZwVpZfl9/4foA7Ud9236cEhbUlZ49Z0/Qvn6Uark
4Kx4nGSKWawjbNA0tGequ0HOiw6SOFR8e5GJpT7AK2JIsveNRwhpOb/EVJvZkT1NpZxwZrxVwVS1
ZBBpjhr7p0LHya+5xKQcukH+2ajF9DgbCJh408oylkdPbZT5PnQIHUAg6HWhRMG4NzCid3+ROa8A
xvYwJcXK7t93FOzfd1mBVgdhqTeaDDz271p2JJb+mfqEhuLmBYoizDdAR8X+aySAzGYzCd6w3CM4
q6C8HUlnTsbqD48YE/GBFciyF2d6vPh2DxUslsjnT+kH7zeScY/B9XNwns81zcysh4ZrQCAq+89v
8iYo5tK+MrzBygQO7kwWoSRToqrmX4JeNxEaDI5QEqRt1pdqHd3I2I2ff5qQVsvyDTihjtBtFe7U
ojTheFXFaeCY+nz9RnTQv7F3uR4naks4HRzzzLr+loKl7NT7FOpaJrrodXQVWI5Nq4It0tfr1QsQ
0tlyKyfoV8MVkytzRFw9BzSq1NVZ9GI5klog+UbLEM7m2WQGWvP4TIC/4F6q6p6ls2OnHV6gDi96
7WnVg4sUPQQXM5ghJEPezHnINvJW8ictagatObO7VR6TUD1ppGuIiaNrMi4pP5BErmAYstKb/qH7
pQ9OtquJ8T43aXwjvING5oUWu1vuSzsknzUhk17MuG8QA6KU2VfCpKXGqKuFM88i53sCsS3bWoiO
Lc1P5EUHAeOGzgs817sr/aaZmXFSSGr+zlQg70Av8RX1aZgw9WtrTTuUzN3OI7JYi/TRyjg9zwjt
pkirxDFL7C+NDBCU0zARdVfSs2kUn279sDRLrs0p44ikLBDopvXK6ntVli3d9Za3JvSiRqWWDjXo
aRca2ND5IMsit4t4XRl0qezUyTq79XPInu3Rxs0vilnLJAON+XmypMyBi7RMtSX9PK6NkeZXNk5d
hz2jB3AeWt5qgRa61sxM8JAGAnKqqcAbUA+QSODYeHMrqcw2HITjzjqCwESBuGujpARuz02jBmVP
ltXu3FMxa7ZT7aTGZBkzk7Z8zm9u2q3KvPFpCLzurKto337aLiJTu+qsUVZFSyMwfdzvYtmB6gMl
aBJ/fRh63iNhlJ4yhECGsQhjuWz5aFqTiYu+a7pH7eCNVQ/C3MkC3uyGWVNOOU9ankqxN4ztPy3X
QoXydQJGyeGHTXrQYm/d1rt62TGNyzCOZ9TJcB65tbYjF2xmEz8px11tCt0U6oLhYCB76iXQHQXx
xyeq+Xrm5x23z0/AEFKwOARqBkBghQpZAkRZL0Ph47kSUkvjA9dSS8nfMymMIRtedLopvPAmjucP
9ROR5Bm4nyYVr+MZ0tOCGC8skiLncYo1u1eLMCPchLyLeYvMGGs+hMo6gulpL4BAkkvTM0wT2eoL
Yl0jtNHXu9JGRFSjdaTf7YjB2uXNYsC33IQT0sO0M/VxmESX08e4K4FppQybgOUF+S+KFTLhOw82
RHXRZAN2N3IwnKxp6AFFn7llzImZ9SzqhsrLF6Um8gwlaxlZOPVT1lpHTG+6lpIDM5umzgxCD+Vh
bLdwlM+6NlqdI6+0ezDC4CW88ot8yhZttMKFv8yg5F21dbNb/1xzBlqEogyPdHvzT8hXfsqeVt9g
NxCE7PWks7i/WocfOZT+TUrBQKLsK9zNEWTHnd9rIG2X2j4DI6TlzQKfPZIuZsnqjR8WN7KK0YD5
RcPrcC+rP0kP9LXKtUVoYraE6KZzBOmd9o9cTlfJeNcNrRF6fLEoDs3lYPCT4+lrI334/fwAXDem
YM0bufinQ1iude1fjZ7oEa1iqyHdHMp9pwEYgXYLP3gSgNCIngHi9pT+aWS4TYwE56y5Vap/2UxN
4MdMGZO4xFJguSh7DPowKVPwDSQ1oTvZZzMlUXyLC/R9713h1liHE7vEmynPClEGj5PUGESsWmwc
QJmdm8O36gWU5NAH2o3xWUly6vXR5CgVHNG3DGrwkH89p14dJi6XaQgI0foP459Xn/gXaRitdg6Z
Woerg9Pj/YNrozuQ1L8x85VSDJ4FDlBs2jbuYEGyObfK6bUO/+RlLYSDNaNoTYBkjCCRsgSPi4Jl
8xZJ7MyiFW98rh4XJu5AR99SVxWwXPEPp3T919AH7U+VJ/MNSk3+LrXZHNgqehX6Yjh8N+4eEGmQ
YOHF75Xw10YMDZBrjT1Den8DbFxu+b5OcnIeqZ7CQ1LoiAf/pY8TSIUB3xhPD+Oa7Rh+WkKE/1lF
WRgXKXLGDfDU0WKI+ea0YGjxOscV6zoXElbyvLWTx/QYcLq2v6bDB6NkwNX2pQe2MNWUO8NJ9dFs
mVRNEze8gVN1HGmaw+hlHVvUJFYQ2ASsNZMD0pRs6ISryf8H3qA00VgvNPCVAK7jRM8i31cDEmJ9
73Sec9iy3wyoyHVimryNieULUAgO52iJtZ4oxsJThI5nkaaT7uHt5TtByWDnMtztJidWE/Pyo2bc
YG7C1cSIy7VGe/fqxubC4vCjsJqiy5IqfhLPcKJZ3JafqsYuiNipnM9mW7TaZ/VS1DVdgrig42Yw
u85FRbj3YgMFS42HXk9Wm8nOx75a9Y7w5qgvYIipMcWLW58/le5nXxzO1E5tPogqdWVIiDSULTcQ
MN2P7LKrggjL51Qcgic4PoI+PVyANi6ukMQKnnVT7Z1eZfAS8NuWaxvG5GzmPm4WY4fKSlRVCQr5
dnFTGfFWoy23iAv7hOQwWga/3D7eNB1EP/WzQkiFz1ANNZNk1DRzuwSMxvzBhivS0n76X9K+4jIb
yaiww8pwN7j6serEanJNG4GTT7bfv58oFAvs6uP6rZj8YOi9XVRmw9YBtaEUzITemzRVJt5KPHU1
ob/cFizmnwgOIB25AB8bISRqhOMu5qXHOX52LxOwOJD3xp7gRM/8wIMvQW5NHmR1V8P0ah2ARQo1
FZ4O4OHvlIz4U9IfnfX4CTgHnW06zdIAqVW+O1Gcg7QkojLaZI9TJFGB8rZhXRTxZj+mkxYVR56n
JICrGZIZ0ynj1LUKaGbhXzU68LCXl8yNfBZJZ9MNaRm2ycWBQF/VEaAJsH8spDgt/3OR1AFVjLHr
JkD7rUXgrODbwbAPlGDuo7UVkohYXp8k/Zwtq8LD9PUhCo9XQTC3pZqZuBpMLOHUiMmKgJDlnBzi
NcZ9vF0dgKqGbSTOZZ0nZKEoFfrBNGmTvgKibsVBb+CsKFe9UeTBDm73IGDv9kigp7Tcl50MqKwW
+7/2MFuT7UZiBVG/bZjlq9fLNd+EWYEfDH1Tp+wcytmc+4EsYE6H2qYPWB/881Ibb6vbsMYSlg2n
UlOBqv9KfDF41eQsde6nETJzHL/fW6hzNVZSThh/ZVql8p90VGQCvtTKRPSTtdG1fhwb5FaA3uX+
FrOI8DyzbqHzhAa5kl2/ws3pelD/J6JlfccZ9QkzKmCMReQ3kF78mWaJjM6DSnwNhLJ2WlHs6npp
IDYQCDiPdq2YSMTmjkTGLGmQr/gkRvS/n59/gmrEn6Mru49uIkHEzFv7M+foPcGSbEOOjwYTlfhh
b3Av2ZHJyrtYSqe8UlMZy9Yw9+3Z60GHdLVHahuTiU02zYeM1ohp8kaD6fvAuS/pf3QHrgZx6V3R
xjUJPGAlvqiQ5rf743agJbH9NwmRTAp3DyX8wuDMlFROyfNpQxyWVCfsVK8Qt296RcM5QN/sEjF2
MQXmDTsvNAxQYdZ7Jlh3wqBEizxN7XCiK7463hee3GAKNo7IQQxiohD1iBNc5879DWFhclhZXcAK
0XNF06rSjci9xAq1sHs5ZD7K2bKA2Dy4PbaYl1kFOGWOEm+dQKSk3yOu0eoBaeL1+k4F3BzgTOqp
ilvwRQ/KsEKH3iRaTlG7WrGpUwgf/jOfZ4gJSgnNXwOntsDZ9HWnmEDYVZb1fZehsyvci/oMqGyp
VmWaHIAtYZ+K1FkE/A5/YluvVHqY/KTKM3xqueHSNfoMh+lE/P+HEnTFdgUYpgH3oXgUcTzThF1c
e6xdtdnQfxpHjEUg74pBCpEyfJIrkCzH7TeYgKJ+QUJgczy01c4gDMVuEdkPohdCqBq92lpO3dr+
vr5cDb7A3bJEmkVjzHNaO43orDz7JioqaW0eeDweNJ3IpKHZL/9onA0anMdVpMwz8Eti+wLv7Stc
1zML7fIOsMD+q6bvlsYIivb92pTgb8ZI9w/D/3g5ESKiQHQPPpSQH/I++9pVFvCH67tCj97RmD/f
UjuWXFX5B6TlFr+4ZxhgobJt8pg7O7Zx3l+u3cpBuNvvvDtNt3se3zPI/51HdKw5kydoMaGQU9Gi
UMdG3c0XTD0Vc3sKX/kWjaeDOEo63NoZIa9zs+qejZeA3UggKkakaf+5wYavQDmXH9i1bRMarP9j
8qd8dcpgLvkvS5jmDKQjZA65ydK8p3G2e1CQHIGOPmJ5s23tJ4MlG+UoRqHt0Nzj4K7bM1JaV8mw
hezge+pthTkqoygwjrqWVdVB94ByBw/2xB12xK5MMCK3ndtXmZld17pZ7bJW3zqLokvwxlB0RhM9
ZJiCjMPIIkzlmC1Wiiw+s0458Xi+UDnP3mqLT/aKnKER3spCRroxCgWyZz1oqLIg8ybq8dOxesoe
V30u3BUVogvVZXnTSIq026zFDkb9WOiApqpTzIuMzYuSDlZTV8bLTEpA1hNkoLSFX90UuNjf1eMf
+SfLDZMg+EBbQuh1ZBqZ5hNCm5/BbXwafEzYWXep9BImCzEmqeAkMqyiy3SOr4MKh1lIAQqV805Y
Ux68vJZszKd1jCq0nMi5YGIcKw8DgZRWHbfUlfO9Vzzf6rclgllg2I44I2os3fkCJtx1NplXIpt3
1V5NdG8hgwagsQIcznS92QH1CNRrKVkhxsRjYUvnfmzKX+7Xp71jfmtd65ov6jR1FPpZsgbCZ4sV
lz/CDGl6wWrUh8k+cM1M2vHZaTsHxxH8rpWBSMEtiLzbGwNmsUboHEsA0FOLDAP5ZGrRQ/wPJb3b
hLkgvuyddEYHNNPEUmKOSODXkL7A53whPiGBA3yuvwTAk04VmskqPr3chkMHqTDMB+fGdpTA/3gq
aZFXAiQE6VB+fPdJ8Pd0W2K5+GObbJJyd5YQZsVBjIr+Z0bjqUnZbqDS55UgwOTZ7UBhRZioEnFF
vPxpEOnhwT3twmh8HUYeZBV3Fpf77uf0UyIS+t9RrioXIxFsgUOlcyeDlK0QIRDC8CNnPkMnQ9EU
Dsi7nNVgAm6pX+w0Y13Eubd8nzaZNW522AmN8NWmWPTQAsMvzlEO6JjQAtw+S4l2lPgqS+1whC5l
N5qOYKUj4wzKYCBPyNS/CFDAIqj9kBPx6hXfD8J/5gl7AhyuGsw+k7r5dWW9Bbtc5jsxoHyI+zuW
W1WSlVC9BpD0y0IrvFw3/YSQW9AFqsVZQ5CpFIyLbE0l3mnLz/xD6qNQzRwDtBgJE+hb7oxLCOHx
VBGAe/jdZmj59s6hJYTa4qc9ceHjSBV2AXhg45Ho0tvojNJVc/2iAr8NH87v7aHrfQ46gxswoA2a
zmg9x8/lKJH1eWSAaW/5T03446dVbWX0lgypURLJtDPfk0a7tFQOn0IBvZcsBXlJ1Jbe3KLEoEl2
bm/RT9K5RU0XSb0ywOG8Ynj76ZZer6XMuVhnERHxNMrXucwqzNcVXJuL/PAALmam7iT0bJ8X/WR4
IQ1uweDxw4APo6q5inmbb3ZRr+LLdRTzSV1xuZJSqRXm6S7DG4PatiC8eXP6rB3UC39YOeGx2g7C
noLAh7HxqmceaOGbHOQiwNvY0zE0xudx9HVzJW7evIWGoK6BmaWm0a1JLWWYnkDH+bhuo48LR4fv
yJ3caVoNQwWuDsgMlw9Wolt/5Hu91Wfgh00kC2k424VZOX5shqOYMUow0Rmyo+E2eKFAmHbPqBpt
xlRlbk3hDqQPyWdqG1VfZHlb0sp4KKWxSRaSS+43DMpY+gGNfLhsQ32cuBZdmc7wyluxKLoJqPH2
jkrDAhOnEvP7jNYQCms8FOiWyafpOYtmnbFzD3orWofNkSy7QLkm8j8XMr+fOdXy1zLZK1cZ9VRh
01FQJscqebtlSXH9Lonq6eReWZVRj8ox0v6L3llt2v1ntl+s2UBAGIfkIxsmw/JvFEMl5Bz9xlek
3O1uflPAkJ+WfHM/XhWgZrw1VLRn+YEzFleS5UxaIyz7Pe8CwF8t1mDZMAsNc+PwH7hsjCA0pDmM
pz+GZW+zaYoucWx5ZdERpunDCps4pPSVte7Uuw2h64dhiaNiv/dxH7tAzHqaJWwHpxPYZntKzdXB
6dP0W3v3L6FeiFMNTug/NJV0Ia25QQztuYaKcCcTGz2PTqhF2k2WBcfVCqmseN5nIehrWQtl4A4O
Tg9uhWPkb8QVsCzwZkW01j7MFjF4+jjAfe6/S9ebe2nLJ7k/zGDx/BLlxbm+qmtuWsuBU0O/QiBS
tq6AUVkdPzZB7CCFRqgAmZ0RMVal2BjFm0vBHwO61susdH5xq9y5jHfLGmaM5Vjm31xISJYhzJQn
LBpA9AR9snDTtyO9IOYyKL8n6Sg8Px49Zc9zsoDyHJk2KdFBWJH5D4Z/nHmX2uIAtedyt6DOT1z3
dhsNOlqtaIilnblAR2TETnDd2ffztqDbpVDgFDyaiC4wXDcakYWu3KiAWDhm58079mO6lRvlt5Lg
UYR8nc2okSG9Y16/PWDknj0wIPJQel4EITRaIjm9PEQ+uyc6RLpu56bVt91tQu971vKrOk0zCFDM
5itMEupoe497SWGC7EIHm5kXVo8gtJy0+Zdxr/otEnVGSqZeRpsSlvNju7F5HRBlsjpuzb0xQ0K1
oPEyVVd19ADoL9vEtSkgXM7ah3ILZ9P1519g7sX8U1p61cfZD4lFc5O1N3CkCXF86DNHKyEZhkAZ
WMJ99cdqRr9esq9qexJe+HiHQDgf/R9OWsAXim6gz9jzXldzBkGGWQFF1zst8HQ6xd7c3I+Vh0z/
R3pNHvOO8vt+u1P0wc8GTAFBs1uiurVHbG4d4m2mv4P2GTusok0wLTfIuNrE4aSVVXLbQRdeMZxh
i5d1tI8Ow6YNoy5V3O6ZnHoRVa1BCuEpP9/lSx7XUlbKEFyjAFMJGAUGkty/Pu74CBLjT+w7Nss+
RqVhIIh8MjS27e9rZHj2OM+CRF/cdqI9fVZQQgnXLrbHzUp7gD7pVviuUB2+Q+hlXCEhAd7dPZCt
ukNn9wqqmDAClcOQ+xgttHlgge36ahVPcxBZHXUQcywMHrXuNnt4Oj8YVrGLJQetwMzmq9aSUtEk
oB/Ckbj5K/v6HMhuHljcgKhOw5961fVWCPpgfiOPlCyZFBzdNeIPRf20Y6vMi8/sjStO6auksNIS
EOsTO5LmNZ47Ju9X/87aXUln+ydWP8e+kpavDwl/RooeTN7nJ54SbSoObEwQfrzE9WKI/t+X5eVC
11UNpG1uNIwSP5xt7xPV+jvmN9TyUgmyhD+ShdNhH2bR+VCGvw8VuzKpn90i6SrUJSNZTRP1YR5W
vfpU7RJfSc8Ixg8jM5xVt4062gqgFcxAV2QwaPqpibURGDaFBuxW5fo2ekk3gIVNUSkel1UohlWP
VruH21OlwvELrUu/a2pLJmAbCjr+CwaZAO3g5LlfTc9Sl5SEOPgQL7spBUO8/kvapuCF+t+WSvr6
vthnp/SaOAxj0+4agQhIF9hWyBrCKNm7GMXh7tuQLF3buVZoCxcijWgN04U8b+uwQjm4MwGoloct
oFTil/d9Nf8LpFIpffsg6uXyJ5q/Zxk/nJ0/LF2jBFLHQI9wBL2KW6Nr6c9Bkjxpw2uLv/FlQVDL
c9t5pBcHCwdbVKsWd8zKLhcgR7JDd9YsBp+bKUzx45uD1gISPDiIvOS+rnMhHoPXlDNDMekrTdO9
YUOmfLiwFuEdZ9F4vSlok130I8VtpZrfdgtDg41G8gqzJyP2wX+Q2YBomXqYtbyuQo0UTdwcIvTU
Do+zhlR1r6qLRvANbI0iQ5fs1vDeBoxpTvXmP32FKSAZucTLf1zYZd/X8aN0nCdjn5BlXmqoI/aq
GjX5GLQWXdrcUSeE0pOfio8q/AZ0fLk6cMdx/dsBRgLgDuKkK0h7cKA9B4kRMqGHKBpfxamJUNSL
eRA7O7ABXUWRYOfgKOn0ood+1SEfxvRYTpiN3u38C7AV9E/7yJ3Rn1TjyIaAFdpYUBeg+OWD1+LX
hg+owqOP699S8on9nOt2WAt3pDr4FrcASjLDtpAfotPaCGt0bW3+4gvAOzfx5bkUMlXfiwyQFGy8
TwPHrYOoEhnKmo5T5U1FTzn4QEb0mES2SFfJY0LQVLGlTFF0In0t2zDMwaFEe81+g8u4olYiNY3u
IYM8RrMoA9MsxEhHMwG3sJfakWalNhKS4nUUMgaIvEZFmW/YuEmuH1BiPdU1uKm/IbVZCJsadg5a
CfilnWbUT9HoTnR4YePNAM36vnDeTlpQVWbhTzc1c0koHTDaWdHFaVuxud3ZUjks1FgEg54Mcc3E
ZlELkB+CBq39si8BvQcpGuIn5eMGo4V2ZF9m6D+OXYzvjxGZWfbd9eYDbVYQ6vDXau8jN4ZfW1u4
QAA/SbzKOnpiKa7J5FkYCOcicDZm1KjosUxVQsnQbRqErUUcqV3hDWyxKB8psweE8SjRjz7oqG/B
W3fnVJBiEGiggcrbHdgVlNZ+/+p8IfiWPKEyLXZlQTdotvAoIcxy2RfmPnv5ouJy1e+yCgjvykkI
KOsHyWJTW6rUPHx2s3c8hKNDVcg8+bjSvFrXXT8jgDC7a2pZyBAiejFdEpxb75O4P79ANm2HEZzL
TirCScLD4qmQuhb0gsPDQUeQcqzJlimxOx7MfvJfy6EcQ2l9cNKCzboTCKscmGL7gU2BQ+0P6/9S
p6SJCQB9sgjhlroClIUyiPPUQbKUl1n6oB0p9TnaG8fDwhydXupGVeHu1avfAwBJ2hNuSKun94xA
tWsSWBnyZUIFf9EuXqhAIET4hOwzXDJOWw8DFZF0xGC9SPUop85fTaZLwVpuSvx4pzbbnBaN/bdl
x8NyTvcMwovPQFRE6zLqR4lIUUA9pv1dcNVGWyC5Lb3xp9A+NkTs1MYr5s8WNzS2aJjq3UTtwTSZ
iuQpoIEcIFKeqTGY4UKOAyZjoHELcwOStaVHx7EBOKhabGq5/yanAp9U0DP93hCcZe5+izXhJPSi
nxm2m4zJjOOYnl9LLY2dA9G30aR45no4+X2A1P6Wt6lxWbMEX14YEL8Hu+Q/xhNRAJF2Wmz+BxWm
IedmBU4J9V65gF75/YL2MuyIeHHeMtstkjUuBs8getaf8kNNbAtWqljER8StNLWYr/wW6lRsn6tN
WBncAGqsG90sCGKKUHLey8lAr+8nZiU2rQbrfJal/qkrQ8eMPSRgs2BSW/s7x72aik82lOQ7DrOQ
HJl9D2LagdTp6vrFaUFRuYD+CcO9K+uhWmGfkPQP54PFwwYA/ray/5jg58jb1nfVaaK6lVHTuXqk
S9FuFhAHD4LhEEzVOWkMl6GnqyX/1bGYCavWC4sIkvLg+8hNTh8J+ciH8w5zZ3Mfeo3EDWmd4Ivi
556RtIM4GQimSloQGrThCCovRqjFczuDCZWJIR683k3Dyuz/1eLv743UTneQwCUVW0+8uyF0XRDq
5Fy80zugqUL9JfaspnMQ0iKoOjxfW0Bu3ATQq8c6094JwNu/U7wqeYBvHd0ZE7lstpRDHIsMBInN
kOPLIQsA7thvJVl8D0r0iThObn8USjusw72LeoNFVpDI1z5rMTxG3zOVcE9C5Nr0nPOKSa2TYCyj
6B/2tWCAOBOUH+gzlJ0jwUVY6wU7+uf+jYtujY9a7RI/jMoGa/nVt6lQ/XDXSXz5oTdFnq5Q4nbx
KHIObQcv1ZTu5iP1su0VyC6wlwnFI2+nYXIDy/KCMMMSNPIIatzhAKXQfte848DLgCcpuRARA76H
GxsIMgFda1bbV4gJ4wSQOvZPUWl8NLV7393lCJ9SelEPN1KiAlR74zqml7cN8w5NfYcMY93J0RLB
va9rzxkxnsn+zpTmcJDRuHKFcDdtdn+61QKsPL2kRQPARvbORYFsQwzT55dSqs9GMHGRSWpB3/J6
Z3JPngfO8haSj7NCWV9v1m3xO5nZLPNrWhSgAKesYnDzbF6zF0fx59NMGlgzQhmsFG3eMwtiyArS
svDafxmbshztq4r+dAsRVNPRsn7VCyyr5LaG5gT7dmXOT3pEh3HZVLQDaxyLhxYxb10RXLH6s6pT
hSnDSouQZspDKdfhmUFUNE/nxLFtuJOFELFexTl+jWMOiNUrjFGT1yhDglhKUp00Jppy1hpqqd3j
ZG4eSa7BzB/OTvYND95ndZohhdgRPIL14zec6ZMmZec1d5jcJ020cgrFP3OZ23n+9tsl4U3UCrVE
2WHcO8NQz2IwOwjGU8PFsRFCfE987cNPd+m0NTSytm7lcY3w4vY49qbTmZ6Po7RKvL9tbsc4o1AG
lZF7UrINJ+pa13xBhVta6oNEPlIs25NkT4Y2jiuez7oTRk+JCpcmhUKKcIOk9JAHsh6m+LkzrGF9
tkTcQGGQiC4KRUnSsJQuET7c8/jl9UJgZ8tfNdPLWtaKjAx6+U7oQlB14Qjy/w54G3qxQqzxiuKP
sGdEsqlD2cGKTwNv2GVQB1RGMwUBNDbNeXZ8VPp89QD/eWdffde2++gsfKFl2kOjHMSofAi8gICM
jn07o+/p1VZiqMqBdHS+TjuSnJ16sslFrY50RuUb20XxY1qWWNH76mSfWBr1yBjyPn2r+6L3TDuv
uT+ylHBRWsPvGc0n295OgKlQk/BA/zLboLadkFNe+pJpm3xlWAFjeYoFpHo1r7bj6h9ePQAJrQsC
mGv34v7d0X5CnUGfdWIfiY1sUzm/jxsXbDxAjMZtcdhzaEjS3xlhquQBxeUYHgwU8CpuH05OJyP6
EElPznagB4VzIbmQIQgpXGHCCu9z4IQ+mimnYx0JjEtPryeAQ0Qc5MKs7XMAuODB9M6WHnG0fW3s
U7tV9koU5U5QheQ+LOCvyoLpX+/F1ycFxWCPZoTMoaG43y4pHf9en4NGYQLbOIGq39PHJJ4GUIKq
Ws8H6w39qHNvQDu33a7E4zCLBHa9vZRqRReRofGUcFw6OH+ToYcsekk1T1TdlDESKUmPmOmTGTkw
Wbcrg3v7dINaN65BNPIAAYB32cyimkxUFAzCWDxdX2aNMU3C7lyMqKtM2Y1zGqn8mQRPJHCSnZRg
0RD7GOgZlfVqn5CLCoL2JGzc8ROqO1RvmuXJmFt/zzy7tosjZ9lKh5RFtntd5b1vWzIr2li92xYm
awrt7PWAOP1ATHNlhE4f/otNAplwOCfSscp5rfy6AfwqjpLVHlPTk/c1iAAsBmF/GyFpp3oDvGME
7CpN6NfvLBOjZXYh2X9YjIVnEUbc+ksupGhrFjlsCqSV6dY18AcJCY0kSES80DP+FB9Qu89btSca
NEf47+BCyWSpaBI4CX1Ed8WyNTvm7fBXcTyfX0MC4ns9ipjtD6tWnwlY7ilZ0Z5Z37odZnQp4Y7m
QPNrznizP94+Az2WyvOwxK6kGFUMyFU/2ELB+GYakkfYUOv77cOd23PI1Ft12IXyChT6tTkGTBnx
6N6aG3y0sUb2tfs81S7gNSheoI5QgXdYzliJumvdRDUkpXPbyuBlWabbhRcN9i82/NWDFrZYZI32
IQ9/VQH6I4dztcRWamVBjxhuA0k7QgYQg44LQRShmuVvx6UlcCNhD89PScZbkrIxGbP3TRRyB20F
Z04ixdR0XpRJeBKzBl/arKUi9e0obDWoT8p0xVpxRY7t3TO4OTpXC38AEWLHNXYGKharOMEnB7AN
zigttgH929zUmxhQ4k+CxYUbLH+nsrwyBIr9AwLE7YRL2VhDy2w/jmTmbSF1kZ713ZYfKZJ76ykp
EbCOhJNoiNzoNRNZ4rx9+TD/24qcw+zNnDrIuzvgdjoi4mc8CMNMo04QeeaW0VZ1wc8Ycqaow8e5
NEIjfZ1YWFB/jXkcfU5AP7eJmtHFLmQVeWy8MbE66loRY5dFnPbSNonyax9iDHjuG8QMJNPXgPad
wh4koP6C1UowYCiRpweUdzxdA2zfKwuyXjfDuNQNCKiWcyfKTjEx94Tkn/PjIXre2R8QOziogbb2
ORWwIkdGnltYcnqC/wxO9nLWNDu3qMLG+UFCXHO3ktcDGPpipk3vrWpe9veicMjAPSlJDtK/ue4q
naaPCLQtKQ6IaCqLH+xIbLqMnUnxwjC5KaKK2XsaYUHrJvkzTAOE/MH42tnRZaqIUQytM+mbA8kX
nEL39wv9zNc0VKfYD27m0ocVB+6LolEgDcklVzGtjxeO/OJAP1Pk60A3yNC6DB86Sa8n8a/D8ppU
oY5vQ4/8mpCC32i+pgwFlJIBRmqeEoHPlkSRqoPD4IFJ2Z2Z/hk78gyB+w/1QSAnpsIcRZDdJTXY
dBmTHFXa0lFWh2xhuWJzZVXZ4j/vXyBLN1ckub6T2JAQVsSMSYZ53GXQTaIglpFB3m5CJ0riR1+K
e++hJCKEYx8NCeHMSUO7C2NtbZZ9h7px8PPUzIK7RAMMK3E0LYKkdM4AJsf0cEFxWDWTJWuc/2AT
2N0/WTcv90khq+DOvcuJJL2IUXB3aKXPNAvmw+ncWahFnVtZHe/L0v7Xh/tr143s9v7XgctATPkQ
w7iMbZgWmIf6G3iGtjV0Qs5uqi2nW+51mhXZqV1IUgTNveaEZChFvbJoBpJAlKbdgzhaVhPaxJbK
FoAcf9wRoRqolyACkY7oIbLDug/YcpBHLilL2b75cSpsvnnKJzxNHmt+tMx8eWGZvqputJLsgFW5
ktoEZTsOrh/8MaS0laZNaILj9DfCjifBN0EaWvPqiun4bCM2mlyGvKo3LbN0SG+FRSJMW3EwGIMp
ZGa81KUFGZ3rxUQq9fkg1DlEzywE3AtXUxE3r/3LLH+F1sdEzgXppr+gom2mJvYWPzZW3qxiVDkw
M6jYGsCj6WMoRFyzjzF28itBFiTadzTgAdfdpCJOosFZKVpL4Bi7IzBCeHPyJgY1IrSruYSrO9PA
frPtttexPpY+LF4vYQ9tgEqS6vMKR1wasktwBa/WrgDafaurkf9zih+PMa6NH1IDXb+vL/6yEdvr
12OavJwWpdEE9BhV2MgzAuaI4kexEIYw+G9Dw65oh7PPQys4Mr0rBVootW91RXlLdb4WR2Fh8ejz
vTyzi1SRcO0ZHKu0jxN73nyQBvQ37fWTyQKk7yo8QNdYO0/asacHLQXzxjlogg6pq59uHAY2JVPc
jSmqm4VfWv1a6wGioIzBnex3V62dwBji654OyDfngJqN7n7Qy7Wu+wHMa2RIAHlyD957JbU05dhC
OCX+oTDiXww9l9fkRyj5L6gI74H75cbDtn98LY43DazStirAluFGg1spSD1hCeBLYEd5C+yrK4Ix
AX+w0rOYUevuU1yP1Zd9IHE0VTn9cJWE8syCsra9bqkDtNgEdZ2qS5dEu8dk1Zv1y/8mtb09jSyX
Y7nX1jtw0sCGWeRnhOni0FVtwg0s1zBnJBPoB7WDWdMD1uQdj3340iXppek+GJ/bMZr9LDbzAkgm
cxGUgXppM692ii/QLwEq6Fk//QI/X4Ts6JChwf1hCT9GAoXT0YoqnzTq8k5zTa+FF3FLniybhSu0
/zz2Z2mFPeTOHmGT+w4+oM4fjggy00DyBVm679cWgwqRtxX0PV90KKnBsBriylO7EmBSp8MxxHNj
CHHm4q1TzG57sQXhlBfQyx9Ib6WFos+SpoLjTxiznTDWkGjqn+8pIVu1cKuWcH88OSlCBhQ3ML35
SOBBpRfGBTPtKlrWac7dYc8lgQlfkqkhVqb+8mSv1gftvsupU6hjpk5IT9qSH6AMSN3tfkqEOCyA
OeZkP4LdH9v8kVFc2MHiT9ymRsNOWfycbmGfTUCgm5cXIjXbkimvlXZtdYSXCyFK+qqVrqavNiCb
LcdOBgjSeSajkvTnyPghMKEBjEea33VadEvcHs4F0oj6ghaRWV4TViV8fWJdBN5tQ0FR9ROLl0X4
DttYJ2WNJFxrH1zO+KQzR2vCtNY53xwbEzo8p8382URIszXNqSLsV4M6XhkjbUP+hOhaiPJ3Ni3j
8q9R84qY1zTrnC7DxyIjNBMP4ykeGLnAA/L3fk4MpcbqJ/3/UpMlH6wg5BPPUisydaKnti3yqdNB
BjUT0NWVwLnHCxhpAohDEdP4BgNFeALBTj+s+zNVi3B/jJBCy1ldyGb43/qW4Fv5pH5N3W0eXDKu
+q3WSVaR4ShHN42bleT+t4OQJXjVRKJB8B5888xbc+hEMzqIIxLZIj7M0L6rKP/7Zk49HP2BNEC/
NA0qsm0jRb8XF89O/73Uhjl0ELoaA0W/6GA67lHrwcwF+ZbzTPDYYcwktYpGUpez0uJhvtBXelNa
RQH9Q57D5TzhzVa4fFIFSnO+JPCIpJ3WJxkR9APewZfiX+GA3quspSib0QazTqWnmSxslmd0Oxqc
8NAHfwupcX83qtqi//YW0xMfa0N2pWX03b16O1xTA3jiLbAgyHuxRdoU5cag+RNUwRsEGB6yTEt2
0idb6VxpAowDeoqO9Gn/p8ntRic16gmmVqEW5T6tGhm36r4NOqbuAyzTVHDwbsy/f4z3Y9eB2Xmm
H/YqRufSn+Vjp+ynaD1QPzM/Vtza3yyNP66dZ+C/qwesYhVUh5tj8jPZ3QOTts/CPLm94iOH5QNF
Sykoe76wUezccCNVfvagCEzxe3LeAbuTYnx88WXn0JxlaoOrmfnJOpivSt7KyibAziyCzAh8YhHv
bbxXyxTw/ABxxHJqSQnqpinh8ab7R9scH5g6ICA8g057kylwshQrCzGz2pdQatRK8OUJ6/esN8D7
uc5KODzbS0/YX9xLMTK9ytB+uGthryuIHUc8k54baQRDh4WXjNVBgWMeUbAE4JWAB9U7p9KGaq5W
RJ+1rJfDNK89q8QcwVf8Qgk9Q6NNTgl4W0jiewcVOv60FAOjLp3DC5VwGYAb68W9OrsF+upiL7lW
kWZErUyqrBM8ggD9JLL4MfCt2LGA32DzdJN4RYPgG9TNoTJqFuKeJMiF7GWtdsk8RwO+RTYKkw2W
RkQtPN56kNU6yi8ov+WsZjwcGwjYBxYyTMVbDKxgXCQXkmOteZqR61BIwlaLY1Wb7kvrxb34vzFR
O81XCTQxrX8cFzHPOnJCzWP44Nga/EFqC1WEyuPOLrzEBvclmqsUOlSPcpsVExvKJBb3tc6tsT+J
uDmrN8Y46feiAeMp+C5W4i+THcI4ukl5rC/CY4j3Fohoq4Ty0pdOsOmenjJgo9xWvDMU8zxYs7Aw
AuvM9Vp58FNKNNV3XF3cHqioHWqMN+jqHo2cnaq2gmGhnDLu6vvsmTK78r1t5n/jbtTlb7s0QOa6
rPyIHORk6ABYHSPCFTHUWFZ9k2KHzTz1M6usFoUNpiMxakUYSU1Adl2xOJPf1DAfDWghbZo/A/2a
V9wu8gYKMyal90XS1x0IaVq9gLpHjn3v32e0bg1u3RX+Utw5mOpE6iqWNDzPge6OgY9/F4OXDppQ
lqn/rs8WrVhIrCmS+bW1w7ZqtmIs6q/TYyBursp8cLN1GtIUbvoBTLjNQRZUweIuMZ7e1YfmyIdO
QLYkiUBG6pVk0RcdifjMy0Zi/Avb3mKaSjbmiutb7zKYINeF6JoeT/2Vpi4HFnJpR+kroe3wH/t5
Yt24fmplB9HdvR9l6Rp+JnlGdjD3X7U4pRJUVJuiSfDDmLwlE8DL/XHTrIvch8Si0EthczmjMLqV
Jj5tlpJcqp7rrsEXLso0yGwG20W2Kk4WwxCSnxf245FI7SawodOfDSvjfEktUY1Jmbzfa6QuSV+Y
zdpRMXwnRPEq2U1LP9/PlyHoptnpiMbXXC7W7NJq39a9lbAFjgtb48r76U35Mi1cwBtg3Qbc2ZZg
W7xAMNI5Wy4Xs33Q+nb0c0GaPSK4D28rPz7k+DmNLFe/c3VEPfEpTNfOampUI7tjNKCRvOr+A6i8
3KbM5C8ZmsLNi8/U4Bi38dLCWG2SgP1YeCmbUH2mcj5smmlvxkJxPpkph7Nbkw6lPeLgek6Pk+Ii
NYbZEe8BfdBk26bNemKqQ/5xeEmQulDvP/rbQhMN5lG3OV4WzdB7bh72i0eSAIQSpzeveEUlnjI6
fFImu/vicWG//39klnTNhCMvslsBwKe7CF0LRpK+HVsQuvJ0CnTGFXZbo7Ba52f1AEG0viG8mPXu
PsWsFdnhfcVkMvyTGRN8HNFl4JLzRmf2VwlBTBMXF963kT61OqNKegOyTg6UoKkzona6pGHIDPwR
vSrkI1A+SLsy0qI9pP73Qiu3e5JgRmZJ53aWrgrMrR/oWd63hB1CowRrULKBMKmlgrDxpIBahRuP
usi7gvhme+Gp4BZQ0+YOIIfsr4HvgCz3WPTrNy4W33yl68VHOpCQyBQIVJvZQyImt/nc3W28bkqg
3j5mlXK1wvc9C6TWSCin20y51yRdxPzUs9xEOuJeieNQ7VnjFfRwQkXRaizJ5Yy5xif3Ht84LCRq
g1h4p1y+DlY7oco14XB7eXREnHRlmScm21+x9HtU8ESG2F9vmbAcoVe5XY1CNhz7QN2egdvruduN
FoLOWM/Jd9ozQZY7Ahfg+0mFQaSGQ0f+6A6NwyTS8m069AX2T1UMoiSQONyuDjFyr3Fbt5c0GArg
fFd5nLVLJPZ4RvhwnimHvYcPW4cFbgsfTUdHov3xCZCVLvPgRknDVlItOPaGgSxTzh3j87D5nj+g
Ufni7HK09OZtvagCOzM5i6xnHOY2Z2PCxeWlo9LIGVT/Wc5aXE+quWCPprWEECmv2rQEDOLMNWcU
6er//4n/oe1r7A6dNmHfCcI3IMDiIpJMuIkRp05J+Iwz4DOCzSO5NJMMQIdIW2vAusWFMQyDjODb
YeS3ZTAUdYldi8O+kSRbjFBPuQo73B6EmCJEqVBcuSGewDjuTEx9EJZUWMqP5/Y/056MMtSm07ef
7+WC+WnxgolrA0hFewzasTo4mrjODp1D2PxKaaR6W9mSiI4cxsfGRcBYHmCNtb2WQZfgv8pia1gp
85E8fVux/sc3MeBV4nZn/LeCP5/R46PKxD5jKvJu9QEakTOGcLgvgZ9M38BHYvFaJQFcA+UJtPwy
28+EQxPHs/PauyG62cp9bQ3k8yreYy1Ev2lHlaSc+5TowGOOY7o+UGZPOuxKMTXjI6RfEZUEovF6
J0LCCPwaqBBdMzxbxKxvEUUNLnLY5sozZM7+XZtntIJDkK7/oN7rgLcGq2eldtOYm/IByJKLk0xL
hgUcULjO/R+/H2Vj+kryQWBrTv2Mu3buaBjIGfh2tuBwD/Cw0A7MN35U2CMhO+bbIgVowEpJysXH
f7r2WXNRmv5Cyg/cvsaxCDvo30lHIgXd9SnSjBDcVrsJ7iqD2gV2+C8iTNZOZmQHA/s6Fwd5s0ue
07VogptQbKdCsNcyViqvSlB9+8ux8gcnCRWJ7YeP8qM9LkW3FeeE2BVhG/CECVYKbEmXUUe2Qnp5
1n4aPpUvxJfphpgz5EJHQezi8mQWUkCjK/OIHsmSNUw0LbGQguPUACHjFvXfCEzFKgBctUmVBA2e
80eXKM21OnjJ3KTHvsY4jtXf3kt62+wupGVnEHAM96pV8INZY3g5ypuRb0hUuOZfFs1kswgTQV/g
VERwlWDl7473ElHW1hqb3o2WPEQbTT5OFNnga5zlrGr1nKZqRpcH8lNmv3dZBJApmgWI4/aw8+NA
EOJbXE1Ij6IlZ1RrdFwFD8c1hf+dLGUBEItPL+AeHkUhsPsCaoZuqZErkR1STq8zp/JJ/ZhaWcSe
C1jGHdxof5pUBJX2jQBUYxYIUyY80I2o9pM+5S6CgiqUjm+KYk6TDfohTnYW8yhFF8U3EUsAGaBg
Q/PA1tx0k3qmdBaB8VlYAwrY0qZriBqufJjYviwlby+DiGoCfavmYi9kgzFt2wa6nejHqNwlDQtW
ZYHzGrJUmBiB06p7HFi4A9wDeMAQ5yrj0FEw2sFWR30dgeBZ1F4Bf5ISQtqfxn7DdrjO2l0CuSJ9
UBmsUqBl0Q0wwhkhZ8So1mHmwBgSu9l9BwYV3O303doDycdnEwtE/ODsLG5cFc9ZJbVdj7r7bo6T
3YGeJAyd6XgJivhgXfQ+CicLb3kAI4QjAD8S1+ooHHUT3WtFNYJP/LmV/12qZ1tpG+Hvoa66N0P4
Bj+Yez01bMxbDRLqGkSv4a63nckX+KCaEO0Uli+LFyBzB57G1byqJhSkyOIBUIvkCHas1Rg3zE24
7zX0YpyavaAE8OU19++VKvfDY4GzeNpkC8tSXJeJkjDaHSXDaPlpwB16eUdC9GL6UFiVnyfL6mS2
oH76uAPeSiFdqArBLLVoBdATMIJ4SF8K3ZVPobtaQjH/fvxZvrQqfYd+vq4jTAveX9WzHKRTHZIf
QP7NSd+7FbiXFk0S0paz9VB6j1OIfL0I0/DymEhcxqYi4eQUfxxtGgHAZnSEE6+OIRZBu0sRBKwi
Qz5/j+Dhorvcbk4SSZ1SoSheSl+GxtWgJCAakdF0wg0+lilYP8/A6nv0yg4uuX0e5XrNSF6s8/Sz
2J3CRI6HWcHbOKbon+cngq0YRd7FA67hQKGgBeihw9MyHzuGh+Ku20fkp5G+xQKdgzOQPjI0HNSh
69K6Axo8cLzElaUXe9YSboclndTb/7IjysapSj72d1TT4JE+fIf4pFXGgAbVBPaY/7kJWd72y4kT
8Wk4rJkFhtMKKUp/JzKu1BvDJnAHtkSWNAFNdL3IT0uLefOaLeRByRASzWt2Gxs1nDQvnBpx59Eq
azNdL58nlLpMu+zmYxv0jDQA0tqiM6aAl/CusZa8ls7/mM6OaMqgFsZAUcWrbtDownDaEW7LYbWE
9n60QIqsRT4xfnhCbHxnpgpL6EloRLUvp/233D6B70TljZIcWfGQi/EY9qubHEH0IkUiUvMfXrvk
8QG0RbAXrCgtAB3Cw0RGNTbAcTWbyyHLp6nRCZzbfa0HJivhBojlVI87n3H94ndXHod3vmGD/ZmB
pNHE364asXVGvgfGGjuItUIb+ApK4c+hqDhX+gJC+sJwxR6Q5zCMZh0mGmOPIFaYgipsptbckV2B
G/vkEOYIKZiyFn1ZzE8l8jLxLyZDkVNUrugbFZP62KKnmD3o7NDS00QB/w+TjIzdzYGEAVEbyAHl
O4NMlbC9Z3yk9VO2UA+uNUzQQWW7w/a8JtNV17m63LPrsTe6DQscEdD6m0i45OraP+anZSoZDNrK
zLWFzanIYdRFHL20+/ME94jR9DAnK/N7KF4rMr36SLNjoZkg0uTCW4VpBjbzY6WYVFl92ulpvP1I
i+cUV6ZJTzdXx4GS4Xt/vKxcPMhIkOiBDWP3CkAlvCxLOCnTABL1nwnDCdE/VEQch8D+NXCcdYYV
2eyYhUSw8Rjw5WHkGTWWd8uuW7vGj5D+w+Gs++VNsDrEV3PZmtLDznfqFQ/4AWdk6mR9NniMv8AX
8u/DFz1jRQrhDaRQ19EQ5hNRyJVWH/QIjt8RG+ikJWzgJz9Zg1H4VS2g2xgG5S+PehRvfcaRS/bI
IFYvQ+Mgs8R8/gcBlH2IhSu/c3EygvSz0Vv7qH4qfMpGiAL07rmflpfdbBJEruxIg4afwmoa10Gn
mGrZL1qFNgVkkn5sVF/qwngpPgTN4nbx6AfqY9ed0toETAw7iL5sN1Owf2ECRQNyrWZyfh7tJrId
W60by8mmwI3Jp3Dka9F09qLWy87PoHbKCZmr4iCTpMnbrHzqKwBMCY2Lr1r6Gt9sZR8GoAptPzDO
VWiKUFqvFpWeKTgcHsYuLM7Bk01IzCRVE30Dt3j0S5/d73HRmfEa9hejCn5NvIwN4pihHuL1we9K
0nvku752tQwEU3n5Q3leaHWBwGUznDzU2cnfv2c7UWKt9kCaJbuZWhVL4hb7CN9oZvBqBHs5Enek
e6uFAWMhqurTpvrroZDuu3gVKFJvAT/JIOMMH6mDkxuFoLeWLHYePFN7dLUC9BrI+rzIkNZ3fwx2
f8s8r0blBE+KSMv106SzkUepaFlNhuOdbQScTQbqgHzfkTRFWRN36CG+WXGozCfRvQEw4eCpvnQC
SwrdzgIYLxfsOSggH14chqkLw9M5yFeDDhLtMeoWBvwslFslhnlA/RJNZgunLQXeAqNxvHe/0YPc
kqXX1s9Ug9Ihx4Blp9OLzp0hhsRjFUaa2MWSsxUM2hVBvhIqTCx9F76F5VCReP416yXoEY2mtBSD
Qf46sv+iiLP+Jm997E9WAaMdkUB0JPEjPU0fNL97rtYWTky0LswvKMuKZ9/E8Yfm0H1UkHhJ9T6g
Yll5a+dMoF1znZ4eH9g7wZ4KxMiYweTkNMZIQAPLkwIK+1RwJMD5MkXrLwYgEgKv+hZ7iWdSCOHb
MTiPKuYOkGkE4K7ngi7AswCMLStR/Grnyj0GWce3rh3oCN9yk9xFm4LLXHy+p/0docFqs2Q+MGnt
S2wJ+f8WAwfrt1GrfrOVwrzfPVDhJ7nOzkXe/LKj4uBSlY9xGjtC+kb3mgFbZ/nfS/plRT26ih5D
cOMXj9Ekp7cr45T4xfkKr45k47HkI/7t0H9n6NWRGvc7vZAXFxz1F8twd41LTxzYU1EmMs0ue104
T3PBuIl/wYEfz1xzYn1wHAitaYr83igKudovCiPjOU5NItc92Y37/1XezmEOMTqYnKiZhbNg7R/K
hkJ9TU2teT7ewLv3tSMyp5Siriaaj8xHDXPKBEfRRVXZZO54Y4VZHzGXEgmzHQAaCYNHWShKLula
R/hvSM9MW6yb/tATSAT1ukEmEa3Ok3Ruz7GHMrGnOpmQIeTHiF2iDt+AyR7u6d2Bk0ZLN/K2td/X
og5wwH+daherKWEeUCzlpRiAXv4rp1g+zCnbIGO289gxe1lbrI8BBgQ+XwkiM07dUVhYtPwH/bWT
+Fh8dDtRXJhFsgZCY54iqvmtuKQifh5UNI/fyDyNfgxeMru2zPd4OHr287DUgWeUldTKwtBTMpaA
atlkoBjUD8qZv3ZKm3qiaIxHApG8ztctCgOuSs1sl7G7b65PnVZ4RzMnpSFFNnhgEQwQpF9Er31U
RtW4FcU3VF3tY+Fhf78WKvWtDHmq3xL2Bn/gzQkPU+EzcZKMrRTLyiZpceGkMrZ11dKupQ7vps+u
DhY9jsiDLkzW4i4ZsTZbAsEoyTfEgsdnNmky3LkGZAlW1QTj6yBc8+d7VtVFdd0eA0DKJCDPMyGf
U7qIOgn3Br+09XAd0IZWpDnmf4KFg/Tr5ZaZmWtLLZxKYfg7vQiV30Xra774d1YrAler5jk9rKrt
L9hdWrV6Q7oFt3BZaSUzNn/v4Ddlkgtuj/FbbS4pK10RgKfjJ0nfzRXoLMjHIsAFbL0PJM5fyW7g
qwux4JOSShung5htfdrDf/LL9PSCKhL35VgDnUgrwon1VqbsJLXFIKIEc5ogkoHRjzMRq6Lm9qYi
VOSKI+VddfEdnYPBuxWiKoCcChxMTXGaX9Ihc88MOclhBpRqgbift1UvL6pH7gJMkBzHpqw6+BWF
Q0Va4M0LwJWmqVXouV3T2WcN6tTDbgoT4NpKDPjN203ldTMDjmIBMLBpdCRL33kZiPMyA0ER0dYX
+cDFFJbs0SCXLP8oEhqydcdL3bQNp7cjuJO8kacSs4ID5n9Dj4EDz9Xe5aGHU92RaRHbtlYvZewl
g5gDxXZZ/klY487cDYBAKX7SdndlIagW/247WMtkWZn4IdsPbrziqxKO7arAe2+A74S9LkVLfHcK
nhkjD89fCSuqXnLAna3IH4f2onsKD6RYj3oWlqwlQQhwlD0nWXD0FEXVgP8Ih8Yp7IllONjYqMw+
H0Ait/8qcgNjZNmpgVLqsKyS+El9ofruLnHXU9poObJ28GQ8ZRCqwMozAuVki5ZbqBnEgeLw7ZjO
xjvL3Ymv8U46qwwBluAdXfBV95a5rXAN2MjsSznPdiUn/IM6pLnPNWA7drS6YktoNCJxu4UfcVbK
//VKzMp49aIqPi3wENngcPZw6oesmAi6AOg/4SYklP+oOjvraUGYDp5sXsHq3oH2bWmJGvQrQocz
cj05eMDS3o9yS7tckA2ErJTXUDrmxA7/bItj0aIEyzvcWuOD7zx1u399TnlqkQ1lGOXbyEzCfXKA
Mvyklb8mEGYqLQCOh1Yo3ecPDVhy0aDA3DboSgqAJpNU/0+K4ZMv0KAEOkCX85Vqz7Umdg6yUYMG
6hySRSML/ZwJNKZnZ0IAp1qdUuDV/Xfgl+mjvF/Qf2cvfuDabOT3Sd/lfWKt3EjI5pSAa4LD0M88
clTCauQxtpefoI9j87XUiwTtcZYehY6UnRh9cHgHzNPTlHHCwjb6bH3HX5O9CvnOr8dp+qqFDiHM
jM0fOCohWcnPfR5F7dbVJpcJYNW9BKSvTgcKN5tWwWwWks56XogjHdToty3hLRydIwnj1nIDlGG8
/zBgWadqy5tDbNI7E1nuYYHZpUAJc74zxb8deEkjJo6jsdA2gn3+LaXh/68SKuDACsT+1WDyhsB/
G7wOA6MJW+boPCChSKEv++qWK/sx0T7Cimn+dWYP7YEs8Ko+akDd4mKY728kuJTkxNn4s4Ft1CO/
6VW5iGAncdaw3PxVZa9Mcz39xhOyVqj4fuGIQA58qgskjb12ieTZnkwtPIiwO65XOOOl6Ea58Nep
X1x/xwuEAJtH8SseOm7xiX3DKNjmJwVcX2xBGElD6DmEY0vGXcRujw7Ynan+JwEVjos+QjaRr/IV
XnRJZq7vedLS971aWUyyW5F8mGPNO2/t9huRjb2guqJ50ZsxwFykjdmWiRd+hFj73aqyeRgcj8Jl
3UVUMnEL9kXrJDU9FkKMs6QPQXDOFoVpMT3R3yzgZFZEdDvC1OXt4tXV7j5sabN5pbaH/tIOaB7F
ebQrNmF8l4ZE8YPmQuvOzyfzwbPHJurakP5GU82QzswaP6XD3VsSoOJWBBE/+t38eD8NV2KySrXF
nL5Okkp10FQbhBF9ccukCgehNZhaS2jgPdwOSmNp9gbZiHZ1qspfWJCtsqQU+pTPnAlpXbcJ4C0v
4R2tBQhjFA0A0HWTQqK0UrubWmI0oGD6pM9qlyy1cdW18gL/K9Y82xwJCC4yQguJH3fzgJrgLy2c
8Cn6tz3jf8Jb1I6kvNNq8Vpgs3/8YoJzJ9R5+dm4Dccf9G7mwUu23KgL94t27RdZ4MzmjWmGZYnk
r+qW1aWGX1ie3fYxzzoMX7D/8pzPjBZhUSXME3D1TRuyaGXb9V0gm/wmerzH86A6fBKRIVLkBczn
uwmI5hr+FrV2Od3itATPPl8qPIXvcXH9s8LNZlFSXRWRQdxfe+XCOd5jaO8QoMA1IVdLkheECNSJ
YaG9WRH1lwE9QRgAKhFA5cTfbNmsINh8CWxwp11nhgB3/KCWNWwxAeI2gCK6dxlDQGHbrg7LJZtC
fRfVljZjEOvwYAJmKW6p8IFEF+gTuJJp2g0hIX3OyfhHmGeyOB71BEAySuUIbe6sRf4eqOgfvyeY
/GaPqGznuln6lZ8QM4rGsDx/jSLYUh2Qy7U065Y6vwNJFwNFuoS1DnKdmuZ351R4Pqycn6NUwwOG
ad8tuMgB9WRRO8QijF7q1QAU1w27B41yqmrBk0MmA4hd193tp6KfkBRzUK94mO2qDZ0mF09BK9mg
tBun8CfBV86UjhIOrTE9M9XBoa6ugnByMMJLSss1PgqxXPiOzAoCfOBxVIzRwoCT4zAW3onik2tE
o+FgbR2lDeLc4HR9VWftXy5W9W3hG2z3lya76nKK1iAFHIdE9iyInlcXHdT9lqSO8VJt4NLSj+2H
ME8yKdPhhz2YY3w0UuAMKDVr0SIcmIey7+q4U8H5nM/6v5Gutfxftur3rdkKxRznm2SpDfezkB9R
qFyjJfCpYGFDT68+P19ulNdLmVc83oEKKFVXqKbwBs/EdqQqT1dUDhvhi5oGurxxvt6SEJYjVwzF
NHrtgOKm4tXVY9QSLbroJucz0pjpCxNxch3ETdecqu3dMW8OxFE0tCVidUEK22d7ynOBeVBWNO/A
ZZOl3iIUxNpdYpNH32gNzm4Nwc7D9lsvIgswwo7UBoP1Kt1x3ND9HaxqMcI65l4hvtOhpSFnh6v0
0e7ZKTgDbtB8po8rxUD9d3eH0knlv+PrL552cOCsogGhsgoQERJFoYyxPyeOiJE2NrnbN9Y8727j
YkEL+LO3l6UwGAYgALQ/TnZL4RpFIDJirNV9r9GVEAuzezQ1+hfj6tSwqb27ErcHV0pOE5b53ELC
7M80u91M+pvcyQxJFRbUQkcfqzCqYatsbiH6rFii2pTdEuupJs0cZuwCLWwyydlOtYZe7eEXEfFM
gb2a8wxrl4DaWv4E1Kb2zuvQUxw/2EeX9Nnn/8re82uQqqqQ2/X3uH57E2aT6BcHPTbDF2NB1IDZ
/OB4atRzRolOzzbb7b+Ycns2txYOF1P1Ywp5XPBQ0BaeacrLUxKHY250ZYM1vkt0qPWik8LA7fim
nJkCjpMAw2aXDjSB5MCqbeOfTBwfqMVhGsg9Uk893p+Af8el3xvfBe3VsVMp/NeV/f1LGnklzQgn
BY/iUtoluYLDGJVRbaMmXTUjSSCdaSCrOSxi+x9YNSydzT/XsUr04QrRwauOj+u4q3i6TZWwjF/H
RomBcM5FKogMJ9RLXvJQkk3Fpk2cpLJIbXhDSh6aTGgB5Wkru5722eKGEmWhcCHeDdtxQPBcUjus
YvibsH849hJxefeY5GkVV4N5ELsL9/LjMxgakj8H8u/QCi2qeFpyvsP64Zn5ZjCxmq55a1Hg5uFU
LE/6rZGJYV8u6G9ypclOqhmSw8+521alCeYkcf/YyHt3qZVSRdRHECxteCDIsZtQb3kFTepjFFmN
1FGhYPb1Nk0uMdGAJFBGV9XW8zyVCFY/t0W1Gcr8yDbBuU+CvXdO5tkKzQDlGeqoBEmuZCJNuEpD
LxaTpXyYCtOaXf2Rnrlyh/B6qdNjk5uKqhjPvk4wn+k4hSji1bkWAqLWJGPtSaCGmvEtkkvnzP+B
jbgy3uNKbQ1gKjQpvi99c0G74R4GN045nn18JMvsdElfhZZF7u9XF7EC/HQ0cvTUc8Ocz8NPaKzj
fjk5LsJ6hvelyw5EFNdkV0A+neIdXLPY/fL9fcWlH8lNU7I2Apg6JVwc8PKcQS4eyYBxDcgouo46
4JF77YXcxIefUvsx4vTMoX7419DY71mjU7k3lPKPOwFkkXdCS5S+TldkCgyk+6a+1iE6jef5STXy
0O47slu3pbq6wo0XZIAzmxlx1aS+qZDbsVYK7NeUlCymj9Kw47j1vkwlA/tGTC/7V/x8L0uCNHry
kZ3wry+R0A/ePSZVMDXeigCPOEMajPcl/IGV54ixFreA9Gl8rMDz4azCRSM8ZSCEno3ov/FC7IkG
Kwo07ip/NIHmrmND1diKpu22wjlpnOpbiRXnE4ZhvjrGcT/gYD5OYTuWEi2vkcSS2YDGcFLHOy0j
kjn3ocQL1wteK8bVf6NLZZVs9SJ2iveu5C346FYnOkgL5h7+l1opkusuSSniLtXseiiaf5hNX30l
IZ203goPhOuEB94/t85pgWHeuY2uGFfSkppDqLKHHzRgnTn+xO/Imd2kfVtiMqWd+yaBE+8HhcTu
tnD+QB0s2NdFBuTli42HgqTzhtHvbtwg17NjyyDXOn43/3unJwbpeWaGs+bS0onM6/QKN6pVulQu
bdYdroYxNAE4Ub6umM4m3gctqksX/7oc20bHTIxzRpFNdzHVoMGN9HvaLbKgbnIEaBSpXhyCR1tm
qE12yFYjatHXCQizpnLlr9+7pjm8XfQ8z4jWYCAu893NRQlENhVfCbAzS9J8Q4yEkUItCSLB/oXN
1c1IWgr1wynT/fD5Dhb/ipUrWBpyuv/ABMSiBW1jaGTptsiGCn2MaSxJxhWuvMf8iyAqMKPCHoi8
pqyduWsli0IanyabMc8+6CpRDPriYdJDK1fFwhIBvhaRGcBvzfwaWb4xGdzFdxj/lhbApUmIOCtS
eB7f1Cuic+rJ6vmo1mAtjdIWb+JiSlrxEFNuG3lbZgm4WISDkga1DnD17P0B1treHBGbHQujWQgV
92fvcz0gU7B4fFSv40g3BciFC2juTBnsndq0+aP95D79lxOrsyPl+krnLi4FXVgPlCwzFPNsGJ/y
P64a5k6ItA5ZQHH6RtsYEpH69mhg5epHrFCzA3V+Zhiu8iGV7EyP/OgNsxZRvRnexDaJsfk0UoU4
NAlUZIBVBZetmIwtfNmhV/BnDkRp7rlF12LDHIm0zhYo44ouJt2q8/QuFRqm9Sup8w5aF1be87BH
mBdaRCzBRjkGWW4SvXP45y69qV3UcSs/tJdZ+hYY1SXkzdmbLYXDPPbgt8a8mfv4Cm04zNSJxzaz
eWanxVd/i9KaAmalP/fPxp/wfBEPhL0UmFwev4bc4NezFit9K1p2LYOWU6feHDvLMuEsyWV6PVwu
4zgYzxXOAhPBYgLGHuhwYICKrAFMCanj9LvaSgBI7sE340HQ/YMTcxX9rchXzyd9FyK02RKe+DJW
JckvUaO3NfcSP/XuFKp7gQTgxQVrg0bXbuW2qQ3kTlhrm3kihszeEDVzvbjLxDgahSXeK9/PEEA5
tNPzYnzK5HB63hRX5NzDCDSk7w4FtLkBoLn8HvVV8Za6h1rZY6SfpRDWx0oA8Dr3Sq1RbZvYWtx4
Cd50BKTpU/EOYN+TYS4qCjAikteMdFa/3A83eQTW2auJig5bMVNWhIpPvZAtgZ/BPp6MJCBMA0aX
452KA+7ZUwKaUCj0Ftf2ZxgOfylqcCXO3gRFCnYgFW9D1a6fSNqrkA7cjhm8LEOS3EXoN3V5gRfR
kRUnVeLPeo/tmR9I9qsEIB5s6I/01IdCy8kaNLwxUnw9eiuw9qhm86J3C9HV30y0TdRZXtRXnHLZ
ws7ovG49StfYEm4PkWd/yNSNV8qpNt69UI7YcZAVegj0lahx6nn5M+8B31aGgd8Y7Xz4YsifVvrN
JqJoHrYU7Lkev1kmiUimNJJO7vRcqlni3mEsQLEnmWZbsflPwCBOtYSKR+aecFEwwLYJUps/HSIa
C9XZGIDDchI7Vf6xE/edPGdmrF7uiYs6uCuF+55aMK60U1++s395aTeRj/5fb0PEezBk60T+Mal0
/KqEL0R2Q6iJxvnBFKSRVg0FQbSreFUCU1s77nnaiS3We22o2wQNUinfTsn2+ZEU0859NPtDd5KJ
ziIb4tHgFoF0L/5pVyJZvPWCGQoBbod1HmbrgpnSmJPgXeq5o2IOV8v7K77J+TB3o8WiOiYhgijV
OJ0NcpUCO+68gi7y9Wi6T5AeWqsRb+f0AvDAGUWnAOxy2ZZQRBxtARq7He0Fa6yllFvSGVkpLXE7
kA0NiCMhOne1fZuJEV39URw3+j0WpZnBeFrF/hRSIAG8FwM7Ss7Efo27U6WekGFi7twyAe8aDSOO
iAHx4TNKpfTlFy6bVrlEYpmUmYDOktToDq8AeMIO9PQ1Kl6SNRqewZvk7kjZVCi39R0qRCEaatPW
BHoFdrzSH38rxF3HKPVIlQnBvl8vJbsNoCE/PoP2pDTAAaF13BrWZNfsBuk9u6u1Lqp6xS0iyPDK
iSw/rV+ppEsAzmfigLStvY0uKG2Q9PObBHf7GrG1f0HmZ07pry9W1Xsh5VHzycb3iHdJvqpx4lkI
FcsJTwCjqyKh3yyEbM7cO1N1+n/x9hQ0FRH17lwclNUo3ofZkUQ0Qa4t53Y9De7Cycl6TJUWmAN7
IDfOlh/EEnQJFZdk4SdFz4As2N7FJmrZi/z1j5D2SdwdjzIr7C39FtGD3RHxs96Kj/JLRu5Cb76r
ihtQaqDR6W8VirifWiu950GuPHq/XVsiq+IKyM0ZA42FoWNltq9nDE51wOWLKJj5hg+bHX5Z0Ein
6rNmXK/PKI8QH/1A8wxx6lyumaVd4KQ+ApjnbDd6Sa7PskEG4Hhpy8rPOEJ1uWhFn/kH6boQrADJ
zABmL8+nTe4cq7ZIZF56rS64/xCbTiYanriH112rMjne6WDDZPd8ugaOk3Uf2Zmi48JmzNHN4bFU
Vg1aY02M4VmrtsjdJbXGfsy8G6ghN4E4ehSq0WA3Oj5E96SohvkHKfvFu2WD/IeV9e6TUU9+/Yru
X5aE8JK9vRTReJ8fX2ty6y2bflszUgd23I+mGEgCeLvsuBfpvJFCDyLKRasNKW1x1arHl3hEY99B
qd+t6bak41vAzlomIkSWpnXClqI5x4cGxzTNqm3u0fNIIuWRiu5qZntmzy1Xmv8LNNkWd2+JKU3E
LyeoNAwmNETAIdUd9kLmUmxExTCJGZbfphoeYLn4y9QTZFstX17Z5x2jelWzuSkIy5OSETV61IXG
4ccfFzpjuFaQ7lE4N8V3mitYkJVbof6Tb7IqfTaiOJp5Q91E+zAvRMRk/8Nc3GskLqpsk+rWGjto
O2Mgb3LcIM5KV/v26/yITtUMoGfZNoorSypZNCov650LmMg/oBgxaH6OpDRbNPY9QoJlnUBHYlvF
yvRvzibvQqinH7gOQVfJ22KM87ChUmS3f9Q+Mt9q6EjnR4eVXkHe2TL5cMaP6o/L7OXgqs1GfCYt
n1p06/uAcF6/crYNRmGsdJD+7pXG8BRsxfXd6/VjOcAVXfTOa2NjoeVDnmE6oR3SXTG2PD5K84HN
cBzRALz3wXvkVQlJJnmG0nPr3pBGkHK19W30U1LZdP47ZPPRQFMpdQXJMnfjSn0ObWKAP4/gn1nG
CHiGKR+vQmZBapB+Ec7CDIDMzE5Bh0aRhOT9Fj4JMufbECEBB/dYzu8KhmEtkhi16iYxsuwjWph1
Eyu84D0DS3w2SUR0xK6cmtDOZq092ejnSN3eBX/nRDctabimrb+q0kZlQm7IvQU3JJfNC3Mt3TS2
SZ6pxjtDzE0lFwhsX50CGFamtOo88Um3gXaI0A4Z8M3f+tAOqi7U/8T4CAKEnTCnalzVy6Q3QHC8
OslGZoZLuy02uxjJVnTdkfTLJ47UpYZwRb8jVE9bNZd3Gyt3MwUEJ2sGxA2rFu+yElkayN2onDzO
DSLhFrHhjF8qdi1Mh5sLWJ1gt3wXwjV4UrYDjDnGY0MOvkrn7X+j15V0jQD1AlDjoPhxc03frkjl
rzoXY8+dCcqxaiZ3hHF5g0CbYxMeBpzrSfg8/evFNNyyXPL2dRgP7ddHok6OIJZ0u1RKRDTNc9bL
vBxrZwjfukg08m2Ou+QqZnE9EMdlRhRn5erby1CiRnixH8Oq5KAZKwdQLgtw7ELF6mntbSIRTZIx
OHTMQDEJSa48eLhNlQ2WftCTXI+Tz2rvsVDNIbu1z6HM+I7jshLVygTAIXGQ77carP7D4yqv5taO
QVrfj/Uwb7beAS5eCR94nE/dSMvnQU8Ggh79fmroStWeDdMc8o8rnCgSS/83bZFumkkngsuu8VhO
HgZyUOwAgQu90jrzwJdpThhV+SZFMeXVTKZvcpS5g2pl3GoE79XSARNL0rouEo7RdaPBwskzpPNR
+ZeKxNOoStgnWC8pkXMS+TJOMw9hHn8ZsYbvCSVrJuLwllWwV2LSsOl/Cc63vmbjgnZo6bzA2dcm
eQdnKuaqFJNyoGqAzUKwfhf2J0Y6WLFfYM9zRvGVucc4gcVFnalSFHsbGHyK09jrmPoOgh/5fDG2
3dl5vr2WuuiVFpNRijJyS/1m0w1OPRMcg+5UA++3+E52lXMaaDBNridtbddGmUB8UdIX2U0siG4a
41SkDAXuhf8HETT42u40e2Yjcn2GQ3+30I5XweHWl9q+PdRnxnnI1RTqIWil5Vl24ZFy9GMpMBOq
h002Mu6907ijai7AYf9rcNeiVCJaZueL4D7+4DXQDBZ2JcH3uFL5Yk8ssLYScIhys6S87lbSigfN
gqyuKrNhDFv4SA4UYJpHG7/LR920/jgFP0NpQAsT9tzhy1NFUwlLUXdsT3p57EtfJ1wty+dikB4l
Vc2TnkL57VK6poicAzreueQZ0A/bxhk252PW/EQQbtrftPUNn9VPAfDJCy42o46QDWu7Ti3DIeDi
9pzKgacJ2SmitB0/7xSJiUmxugvtXoEkM1CDTyY/JpTxRizXoX0JbT6KbiOhHJQwpbxwt2sWnIX8
OeJHCSz/pGCg/3gIb6QN59pHrkIoIkRFp0pGS+YNgTLCYu46v2NHKw7n5o8FwQxWKn6QAkS+MAkt
7CLJ7OcmczwWkkcLXvb2KWhM2EOWGbKyg5AfPT81hADLFVjdrYBMhryDM8TKnPpVK4BfMqTFnzSO
staS2Rkqs/x/C9FgHD5XYLMqOpBTQIRu4O3Liz5qrw75fw7Owlq6JM2x5sgqVKZfo6/jx5S+78Ij
1lbJ18+w8xg+337TLbxAPi+mvFROJMLQNXDuaCiMYyo2CDKfGRYpWlI7Aaz2g6kJuOOHxL1WgS/g
69I9Mx9MP7NPEmTq4h2zZyw3dLcn4WbRVF7spty+nyBYblyyglcyR/q8ejm+rFCFTPROwgQhoTaG
x/1qSYCXxpOP9k+ArYVhWuTKCbVkBRcq/OXVhs4HcuobePO1wI3eskXrzqK6yz9rkn5/4EOfKe1n
0CmSHROlfmyCyunS3g+eFM+7Q1WG54sMdWlm9cwQKPDxr9tp1fdgWQxpWkmXGOyIlXJyy8eEn6VJ
3ovweEzOjx4/ATPuWJiQ2A5YV8fMEaLvVv8og3CgJe47oWGqpV2xcnx1wy8prH6mdX2OO9skLy7t
OzqlWRHETu7X0TKN59s1kOR+k2/3arowk8fDXmfswkbWEKiMo7u7QOTuSM5FU2360zN91AeQ3ng6
oIftOv9ymG8aX0Nh9w41hjlhM8683NQf45qv6YBBm5vXLI3jBmaTmJM+OraynFBKRJ+A6+IfTwTH
lCx0kwwW8lEweVkeqRSIWet5ngOp4sXSxlW8daDtXl2ntmg8onRPfGGrBn7rqFoMGeHX8SabSFuA
hChTkp+rifR493r2/YfBf/aouQXGdfjqSWc1io4Mlwh+7fV+mLXmkX+5Sp3+I8lcSgFz31Hrz+I/
uSr3ai1NVCyVw/TlfXkVOGRkmjk/ioFLAi1EIDXqRHx3b3iS7HoEuly950ntA4xAgEUjd7e4THkb
8k1D/4y20ZORaDSIkotZkbfrICZrKj1sbODmbAQceVVXnJ8Fq5V26s2AfkN4KrLKRR4Cm0JG0oj8
t6R0ZKXt0FLhcayqYH+NauPAySnOikHsOepg/+JYRPsAG8hEb8Pq1aYl9yZ4jmAi0F30XQ7KY4Gx
y6UqyUFdBPuIL3Di/q4RFoodDlGq//RXSvQvYNvue1l2qi//6Wa+asSYLHmfIYsNFtAX9zzIBd5G
SRbSklgsMZnt9wZgL+XFcoF/o0DKQ+wgMASaed3RwI2Sd6v8IkbHiefC9dEOYqm93ckTqlouAdq4
mQoDlzoQIz14cF9yoWXkANO0Nb9IcfffjZTkJFJo6RIohvsGgSqD94L40PKUZDmFK4O7h9FhfdXz
Q9R/Tw5hJ2ELyV/1m9WfBNhlUluhW/Oc7I3CshgoBU3bHhA357lCxm4nXCtk+EGO5J+zp0TTjwww
7FSt0jf5zpaqzenDS82DxAdHcXTL1vm/9f3eio3Oxr/Lz4yf0AyKldSjFIjLabrwlgGKBhMg4Xji
BqFryuD4uG+4rpK7Vk8lpKNosvygpZEM6ODvo01g6wBeSTPFE0ue7MYvv0w2TeHz9gt29onLKsS2
Qp6yZUzZmomYLvOmIXEjQk6XbPehfiwd+kzyQIN71MXPwjaIMsBL6dfhMTsXyHlmBIg1BcphqMeR
wFnpm0rlttBm2vaf0NApRC9oUEH9jE77gPyp7HtXAai5eHss6qH/hO24VkS4eJqPZtfAT83kP66M
uh0oSbMhHkPRn5lUC34McLUxNMxyqT/Z661HqAQv6drNJsNwI6aBTfC/Q4l7KUrPA85yc4Pv1DRm
tGdThMEluWCD+4FP/LrWBCTj53X6JN57lBG+9tT1dhpSc1Oez04UaHrstepYqrNbHjKiJlQ1wAjj
B1Lx+71jMAWSBo8vOszl7cLyW3XMcgOEN2Mf0MeYouJV5TsPeoisytEL6ljn6YoaNmrQkVwWvJeC
0UgyHErLKIfjVHS00NeMpO8kuyMRl/FYYbCUeyv1xJnILbdh+6pD8OUenKzcjLm6S8uN1ZK5QbQx
AWA6RKR3eoRnfI4sYOIBTI37dmr1oK62voVKjgPwgf0OhSZ/eYAvvrdPYSzMBJt0/srTXmdIAG7/
jv8kI0+czoMx2t8HCHzygc3zLKWRLm0KQ+nt8oN4f4IfSA9i+eP/Tfhs5NO2lcEfmhYunHmgI0IO
Np/wOu1euiFTJAconQEOBiyhh9OuL6X0CpJl0s0D4v/GmEQOloC25sEBexwCHGXimRG/CSV+SFZb
docQkLa7VWDqGl7j7wP1YV6sNDyiXGPXr8gORg18GerYosMhQfbNrfCCgSTMp2b9AhXcIY8+/DJV
qKez01mvuAsf5CZxJz+oKoN8xyExHM6rfDrUtpwtMD5IkgIzR4O9S6RmDdss1Wx0DtcD2HUmkOPh
LEYrQ24CshXsqjc8S/4ChihcYHztsfnxLmh7JEM1pXf2pQ0FzpnuZ5j+a9171wBxfshLLp1bgbwD
3IxaOO/QJ2j6YDb7/FKeeXYqxyQi2+GWMcmSwKEyFoWufAKFRxlkVGhHoHskq8rnF/ay7IcuTxBo
msC21ai5xLUqZ6eE7TnhgIJhQVOXmzqWYcxYtbZqheFC0wINGFgGhhcd93U2QVzLXwZWauwRUbFw
lHdtZojGPp1PY8hIxpfK9W8Zhd+gbXmHzKopC67GTMXfIEzpBwUPthtaaIwyL40F6HI/mmRe4/Qc
RDYsCS/wjFRbIjC9ccSZVzoTLZa2vYNzFYz+Iw2sMy67acSRvsIN/mqu2nfPc/O9gQHvTR6qZeO8
oRK+Htub1TkMdMLAUgb2UGHqiwJiEt0NPtMDcpKxJb1vLiOccCGkiGPVmCQ719+cwfmpxiRU+4iO
XR/u/GzoR8ZuBz4ZjS0LHKt3rg/KGgVOzIpSMJKEapkxabT7oDvqzqUTCcQS4akNslG13dyhtCNG
xikTXFBhJXX36jqorvf75yne+zvAvXUUm23QELmIK0co2yScoAjeDULvZcDwQVXaeWcKyMiIiP5D
zWDoRvr61iNnW47mPBsqHXMoy1SGXPUj+aYrR0dcQLt1hBqzDDVlVz9AvN8ddEUIuJiXqgQZyP0S
MJrUpKa4rHXlUN+IiWGni7jWU8kv+RGsayHkAFiiZ/JW+BnO75FSYkVBjQJA6thuGxHRWuOseBB1
qoRqYbvYqhAttYimZ5rYdIs3UEAg9YRznazuuhy9COfeyBpMbFsYpBqef2ByyGyBsM8995pd7UHv
CqAJXVtvBwgOEEwfdSDxgJz3plsfNLPmU7PJWmYSjs/YHwq28FhywVG7oFqAq7kMpYxB1zFxxIwe
Hdq4fQSf8HEjuZ7fkwfxz1mYNfxqBoMKS3v38DaQTdGuM5vtrSKhHimxZ+3RbZXQ+Voch8Lhlf0l
jO1eN+zN2je/c8Amf5BjkwcsM+4MQJpTmzQpqDLt4nTyv2yHCYykvK/rIEymf1toc1Wt7TiKAwwj
vDQkXRaXlI2ceF2gBavM4twumAk7PFG12LaLBn6idY8kCpzHaD6GCb7JbkdO0D7Ha5bJSgoheGSr
BywY9IL7rZhRFcquAZP0sIJFEwKgbTUIREedyfUV99Vp2ZUClVdBYCgFiFbRsEBwZSGFm2Ww4vnm
PwtsR5j125il6wgiwXdQ90AsicBM7FFymb5uy0wBnHJvDiP/jmuOCZjcLKPQ1lymhz84i4wV1ZXW
0i1ikvu+GLaMajzvkoQrZQjRc2SHZvVPLpjbWzXq97lwGU63Xn79VC9GMiYTy7D8d4WIkbhdgMbr
HueSJCPLWWJ9Fkh2OrMokx+eFUl6nCQ8H/pm7IVvy0uP0choPTKaa8KyQw+5WNO4UkSEnLjJHb1Y
rD2KSWcA5w+k7voEKXlmkxRFCBd1bYm0M9iPwWZxE2I3RZ1i0P6VZvLm4BBncn0So91FM5ErxFNd
pnolVc4rbTk3KDk6rPU9jwvYGUl5TS4N+Z5r9cEMDgwG1E/PNZpNd1pjQyaYrxQ83I/Zi1EfuqJ7
ypt5bLSWNM6DGGql0Z4PiKYiwKKHd5S/FeM3lQ5+ckFW9ZuoItXDsUrWmQPHkDvR1+bqHq4KUGw4
FhXWIb9r8jPuYpMuXzvthg2N7MSyYge3G89DZ64bUkRnjNcV2WWs1WN6NXpfMw4RiLP54MIi/Pjh
tTr67bbh04jCtahnibRlSrvGuAfkRbYKdJdHn/LaKmR4svmkHPkTKLBkvOUBgg1aj0GS3O/Vh8xy
4H79jnRfZVESyyDv5wlvrESq6y0lTMSxcnCe2Y25oDE4cU70e/46jp5UmXhsjckurwb8bXBaFWsE
PJkan0+FCW2pSzqFaQk2TxmV2KIrwe/hAuongT2867cjK8thWG6EUOdiAfjm9PQJ0l0Y2fkY1O0e
l9t91n3wvS5pqIM10PMbAoKzrZn0fDu/W5yBMFp8SaCrjNbSkdBbQfz7lvHQKA9SetfJxVD7Tfex
kZh3BC1O7jkHgXVVF6nLBhdOLpUKyyVMPONdAN0eBx1fyiZ0Qhx21ljw5NBFtzvnwQFIC8NMRJ5K
XpeKZPJXWS0CQQepdzLJl6T4aMqUKl1FPGZfiK7D1u33phKe0aHfCsLCuklqaVS4x0+ktlJ1hrbJ
lsZbN7g9dw2eBnZ/AVXhvPSn4ZPymTGPRNP6FgIS5QCLIb4WmuoOs8YxBoPjD+JvnWWSG+3id138
UfUOvWgA02Vll87zx9PZJLasxx4QNBNb16HZPC9xiri0uVZqEDAW0d65fNov8tU4Ey+zTxJyrxsB
A7h2ukdeHJMSsYzuXVKFQJz0wHaOqv/KyNUdOL1HRFfZjmnooodBNdfOCA34cIdvD8PDDeTz33/B
7Q3F0KZ215nqTWNqFuokr1NN+CgmMAfxec2ERB1MUMrb0x6Z2t1iE31FXX0WtyZucZeyRb1eiTNo
c9rHxzrbv29mwCZnNL3zvDHcwCaldw76wq4kG1MBj30F+8IQT6h3y2hTbiubS9h1BS6Cb9dE18Ff
lCnhuTjm/FPBogJWo81CPhblg9EFckj+ZINdwDNHNVKXd1vp2limfg690kdz0Nt1FIkbJU97xOys
Jm7JrAMgo+TxqW5rGnENA9KoUTsITZBvWOFGNoPGdOPO1UHOFangUiLQcW1AyC/mSAdq3J15j9eO
6k1fIOXumZn9aFjhtKPW6Nu8+dLOe7YiBwI+0qNcQCoPdwlqCU20rZG7CfT0Y8HBbEqoiZQrSYP5
iCvBgUHfHpJpr3A6i2usYMlNYigG7Vxp9BlBePR6ymq/IxuXx+6UZHcfwpGSC8BdStYxro+MdDgG
s47pMwi/dS4B5CRpmHTZYOx6QUr5nrUIcguTpnYYEgKarHOooOfZexyB/felUggGnbGqImDJomvF
KKEnNFtsjcPEKXs7I00LLIXCNirpr0RHd2+JsHubCq+MOkDr8TmpIRIHe5ds70jkvt/I6EujG8Do
5riYhuTSmKn21l0COaq/CCjdGvn9yMr91qO6Cxe7fvQw87Iyf3udAtMTJRNvylqvNDaOY9VpDdUB
lt048JwSzeMzq9sNdfJ/F5cpBHdp4DOTXxTo8QplCEDOvxn6MoQToGwcLIEYtl/px2AF4KZzDtLb
os9I8x5pZdOiTQiuqjsG+ablwyNLg+LrKw9HkXQ/m4JgBuKztczfFHpdBOICMMxfd/HUV2AlZXr5
LBsUe5Qs1mTikPmV7ZmD1gZmCUIow7eJ1SJBVlnkpX7uPEkeVZyGj7+eZbQjaquTw6GjwId3O8YL
1SI4bQQfFDOjoH/04dZKuWGCiOFwCbL5bEquZ9p8Juy3vLGP8HiTrzEEaLtLBc1SYbC8vWHD7ifX
dU8W0LIAqRFGEMHBa/G2PHajnITverbjzYBglDtgLddLNjioyVcYs+dWhllJ5WnkaI6W8zUjKD81
olalqq14SNjGCfhd/8kz/9bUsG9jElRDeEJ7IuyZUHy1XUlf8bLrZYYFwTonD4FGRtCKP9Yg6fbu
hQB3Vwq1XwZuTuaQn3nnshMkqNLP5LQgg0STrUttfCoTY6Q9xwTdrhjT/m7CKrpCwYDUWlEYD5hd
yXtcdOclem7yt3JvugdYQc0JCpErly6Umo08uG6fi0mLAfCoikBf7/s/9y5/YSEauil+ptSf5gVp
CucWVh0P6qGPTHAgwxCJtxrwxvPRwdzx6AiLko5J8sSC1sK/3aJNr7/F4dY8aprFZnpY/aZWY+CG
6iL2mZgOZDe0N7YsBudMacsl08dne5MX0GSTpijrTqgCm8wkTxYxe4iH5mbB0mC2FbUmn32N9WcK
l4mBNXXV9+y+TWO59EpSK8BHWDv2wDP6oMnkWDIv0okf0xoZS9kYlYoBUFyIK7yO/+7JV1klg1Mu
L8DJ+/R+Np0a3rHQD0yuhgMisiH+WHjSdIusfHjxE5FdzV71lUEJMs8XIPPCKC4rMA85/RacnZ/W
zJCcp5WqJCPHNukQfQidnasKYthcPbmlDj4oxpLJsdUpVeW1UtRivkbscbt8Q0NFPvdwVmhN5qKm
N47flu4uVz0mNUBWSRWuJe8XHn4g09FHneBg3yuiMxBTJwAT2ORzqI75CwvRADQe1HWac4N7irSw
EVE9igKvW/VCEoc0ypB/ZeXXR9lSvNWxqFm9vALbNp8vUCcx/05VApBtrxEbInpSb2zBH78KGKEo
IyI+kRHZeyqEVUSneBZXHa3Z0JjLRBPKHeiGMaCvlsq4jKdUfRHBJIM5w4Kfgj4/9I+dgF0cmLBo
f+ztQRKweQ0laiouBsKZmfxRk39JFGJqq8i5Db+b/HdO/IZqHTUuXyC1P2X8M7iIIlTLLPx/bUYN
0U+ZYu8UhUQijo8mwv0HwpvtXVM4oV/tAM2GA9t4XoNor5SZR974Bdonlp6nUslKNfns5xkTknJB
SiszkpSnGDgPmErMwXhGEDqHX+tqbN9TMA2hif1auGU2TisLLOm/PyzWtFTwrOu8y83WBQb4mBl2
3c0vAyyt1if5c5I2eaR38YTU1EaUPFuRTKTQtH/GIc/6CPwcV+suhH4FsJ7u2KQSOK5025vh1crD
l7Xj8Qxmw9M4hB97eEjrCB18AmTR5D6XDvyj2xaVHCdfGyGYh4gSzPbUrqh2A3ITTadHoRV82hIC
vLRn7zf7WJYICwgtLeBLf1PACM89kmlD4Ny0D4pf0sYY6mdl3bvxXBDZOzLEvaz//VcfLPuC9JUF
9URhD2Li6/fRztHxH79RvaC+SlOD4a5HtNzCi2HDpQgCKpqtMEvsNau5NY6CHy/K21hj4JbPC0uX
XhOuWkQjMCEpMrCAUmjRidHK2C6z7P2OmOMi92VQOOOceBUgjncnQjPQ8N+kjr6O+hB9sgDq8zCD
TQNpumYANlU8t0lI6AQ3HQbyHXgpW7uOAJmWddoGtJF/r7jyn6X0HyOuyRIm14z11U/RgA4iHM5S
tQvTxksyrzIbiGzXBGUZPZyeKXQP/1D+dhlcZJYkG6oszFfwbBa6zkvTXhbXhqlVB4vp8gJq1BjS
fMeofTyhSgQutQEqSLlxfpN/DmUxRiCX8yuukI7M61/4mWizS2uPdgJiaHUa0YyoPCif8Sphe84h
WZoqNqd+AtpAb5b6C4VYbWok1V4HKajFUSDZkpoGBTvw4593Qlivj+Y486R5OOuulaq2e3heQ8U2
zcubr7CP1RlmrQlWGAH976s3rm2dYIuayCViqPYE898M0+iDuRSi8e2ZFaeKElv5DiycbhODUnAz
Q8MYBTjRU+E3SgpNdxUYLSFmj9Xd/+Qz+pZbl7I5QW5fFHFXhbsvLguh+r0hn2tMz93CbD+eYdXe
rm9sX5emlaknFT0YzBL8vwRfACAqcL6oxlg6JH9YtFQZKiWtlcNtGg4NAfB1bxXYimZHKuV2EELV
kVFFLimqq7VjqG5Fzi60njokoFuuS3q/TOvpRq48BfzYJHLJ5hF7xWzsece/BGmpTpbo2pGttcSm
KWby7AUDPN3zmNwfq1sxu2JPFNBr5kaiwHcm0vG8XnwnxFdy94BCD5CDSAQ2M2Yj7JOvgf99JzaA
0FZIknxLLC7kroJf7KLbGQw0c927c37sdMMfBP1AeCzcAYhr2iUhVxheua7NiyGYXdQhpixKlh0R
aGLSbpMk7Kza1vhvyrRAs9kUTneJ1W0saKoCGsjQZ5vZxEoVvzmRgBPf1qLdrq8V5gpoYXZJo3LB
0SE/rM0kFDXGSeZWFIkldH08tNUnqu2Ac+bZDe6IcqBsZfMh6Tg1S5w29ujW0dLywHQOa0GKv+d4
6nMWKyM631SLhc2ILL84bYgdmkEx837ps6E8nLPAwrciET2maofHegDnrICY86Yh9HDGcGkGmAis
G0cD0Cc/0A2gX6LsV2YRFjHK7vp3oQfPIMB0ad/j4DdCUx4lrHQMuxgWXOmr5GkK55xUnY1Wneax
DepMdgFP+JnOWcylxbP8hEfAi3voUSRFkqDCUqFsorpwU4Ym8oLyMVgkW4TxdPluhHxw1b67oUT5
KquvWbLEzAlhvjBA3QEY1gflT+JLZrALQmNT51lQsg6sTDjQbSVSSJKxAPweEJSURpZ6tnL0+idN
ub0IhNpxVkTMG5SMPE2PxvNDsbgRenzZOk5fkT9f7X9vTPhD6G/iR0Z2oLzhz3V+85SNlAQBb1uS
4xMZz932DaDsINlqKHVstF5FqLChIYN5f3gXNHRFiVhTvuElGlriY2cwWBFuf6w/rK0ZVpAZUIGu
CISKBgFoL2wt4dJAme1KSSChYhLTUyB/WLhfIe/k3KTdjPiKxBorBERza8Wa2VdTQZc5PXRJvjjg
idTn8CTKHAcQ5QjaWGJK0SY/hQVPSvfmbMd1UQZQosTjIXMR3ne+zslmFPZ8Jiubw0qVBC7fLr0m
zavCboq/rqAk/A1rUHB0a41CMVLmrMGGTU9OpbAWOgq9F7X9U0BtGKo5RimS8gNOSFy7eQQ7A0I0
0dEw6Vn6SM1QBZRq8IGN0H95Wt2YTxcsMnB+/v1vOYiH5X+BSA9Vs4dGAhHndGtY2XjwWAHd4YeZ
tF8hN2RVy7NRPiKjSzkgO9F5ahFViPIFxdFjF+ZvoZ0ga7U+ndKJQKXtlsO/D7tCbqQEcQW64UhW
lBv6Myn9tvuyIwQYmxeLQZFXiOP4e+2gxWa1xPSp/iT4LZKvcFESMSl1NRB9RKqw+YroVb7Ivo2f
xEeRdz29NaOBs4aqzQ9VQB9sZKC8KceNBV7uxpvukbm+KlffZBTzTsTxlLdw7y0CUVsMLbSWyoAh
nqmmUaqNTb9vX02MOGfOJbKNzJxMU6q3FLV+p3Y/KlARDafubi0NPdcuhxUty8si8U4K1nFiq2bN
fZNuptQfpZ+SM/mDEU3//epmiONVbXC627kYhZE3GuxEAhXhVdP0f7wKwGqY5Qdw27Rk9W13TNMU
nz6gnGbaOVEfz5uc03msSnkXDADocYsQZ5x1GaBs+iDTV1/Zk5NheTsialsv0Fc53B2afLz6eTcs
SNkFXsIUAxdi+IWVcUnHC9J7nPyUb0CsLz7RkXH9nRw4GQ+mCDu7O8ZljGg9Z25ANwMz6cqPOXtu
V/zIwim+HThVT2ct59ZLwAq75eQp8aJE4i/F6IFDNjTZXiY7/LsLHNYH+OAtveeW3kL1rls+jSNk
3At4yx1WkZM0jI5Q15RQsj4wV/qm9w9nnSr4Ndmw6p+rzUKin/FnuyaWOMHCatGjgcRMy6Q+e7Mp
WBAb3o+wASrVGFf+17DwA4RtHO+lvmvkyvURRbNc8qOBgfoFUYLPJChPuvUJp5v6P5C5D/9IwDta
GEWs6LNuwsj3LpF3aHsKVUirXsB/TtwoLUfRUW+jvJNuVTqMQTp5jROhlg+gizQ5vUqvZkAyjudO
Q46fUos2DVeaCY0UafepIGHsWzjnSgAPFzQoZWP7reCPnICAoqopt5YrY6tHfRDWzR5+kJXCWyLv
8rzr7K6I5zxNVO8encS9lp5SnMxqt64mIzwXo6xIFCKYNHARDRmhO/ybbyMTwOe/8xrPSgBtOE74
n1yfx5bLAlontPhklUwz7SoJXcYRAPNVQxTKFetcm3brazdTxfBuRoP9xwTZrI4zP1J/ENj2WyMO
KuN9ig1D8xf78jMR0FYyvEmJRUY6B/U4XCOXlbhBAdlV9iT268nJJ7YttQX4+BhKRvKXxXw7AOQz
l/cULdIT0NK2g5Y6UeEyfCqC9ENk6yIdJOUSjqAAXLnmkOOJzjlCLv0LBYBOOsrkMbnrHNXdpPvE
xDKoggSy6ywjPvXjREYCWc2jte+bcGFvEgPVUdOCzJQT5ww1L664b4vKeI3vfshWMQ+7m9UZWTg6
jj88o07s3IXSKbcdqkM0yQKa3MXCJIudzTwOVsi0Xlm0Dy3Jef/5XOq/2YmUJomfp0xZkqWm5ldA
aYcKNCvJO8DRM/W9pOsRcLZeq7gPznPBdtNwFgCJzjG252q2OJKeqRrParrGTuzitLBLP/45W0rL
2doQ240UZR15hiU7yJspleUgIRtpBWJH1pcE9tv2UIxcgw2dEGTMsHsSe9whZS8n6ZbVEZuMKEup
cl32K4EqS+6wNCnXQ0V7UUWP7Xys5+rcXflM4xkDdeVKTiGVHkmxHyy/nS9XOsOEVcBMinFhTa8k
JvBMgi9JC+O4T+bA0fipR1wtJSln/HhXl5AFFY8upJP0i4LIwUiL8uMSlU6bM36lybMxJoJUw2jP
cQKNF6RecYMucM6OD7q0v0QELhtseLJXzqNsCW5PuGDVdoQMkBTNGAmkWn/Mi+ywksfDJFnReUPC
ZS8Wf3tdq35J7gzAe//ecX+u+O437V/+FHJkxHemojS0H3wbrpYUiJEF15gDzU69NSPJ0csmjGBy
hZpw1JRe7iS88c8alFLcIUAz9wpiKCJMrlirpxk9UnuSk3NuqcKZ9NxmjoC1jinsqYFQFgxbJYDp
Ar3kJDbHLM5c9iIgmbf+j1+tC+WXfjO3pMLKoLF1sXG6EjksMmx/wGJsrtBLdkBPUxzH7XvVE4X7
dEZJvHASV2SmLH0A3H/ndY4Fk1tc2j/9SsH8FrcK1JvvJlayhPFwVEwYcagMaPDfcKl/VjWjnQ5o
2xcX+kYz1SYIUaGRd/L+OM+5uGnCSxb+oYfG9ihBWkwW6EcsDNkywFKEhR4mtWg2IC/+DLnzZRG9
eZtEkRresJnDjbS50dWG/x+u6p8Ss8/LVhB84UYuRdSt/9qaNihDYhfnKIIvl6AZkoH3ia3SB+RP
AAn8l4QCxRwQi06/+KbmAltAaM85ghSN9msa9pC3ygX+I5b/qsvgh8JXitR24GG5dq1LYBmvvzjQ
5GkIQjxge1c+VuCg38gAADttb6iHzqBQG2BOVkSjqMENfLT5QF1fE6AtipKX3migyJqF7oXB3sHw
2Vdimnv6qTDIZsehPvy4bTrbNt/ZdEGhs77/EVdIc2T6i22snT0W43QVCbH7RAS7pFu2c4IVlfM6
EwZ9w3bt1D13z7gNkRgXZzRDHI1NdHYCveKa06E29tD3nN15JvaRaEcjpX7dCfGsCYUGUCNcrHrz
ngprOm1kSugyFfYyNejHLPc9dTE/g9lkoN3Ux5dg95Za70+P5Txu/W5GFg8lp34m+9UJHc280ODX
2D86/Yeiz05Y45I3v1wHexvjKQWKDReWHxDsqpRtWr0hCZD0lLsn0J1AJg3XaN635/OROSm46ZTw
1tdPA8BudLN0xkAWYrMDe0PlfawQxDyhZxZteLtUagNZzChyy/3GLQNSLRb5aZKlZk3/YlxEcQEK
GhwjJWVT6swus99sgG1zvBEmMCPP6ru5BCzr4dFe2Gq0rJ7+356JWNP+zET9RvgRR7BMrarIBfPT
XJnd/qYyKUK4N9u7fs+QejrNrmUfM0/runP2z0nz/4kfNy4FjlYRqro99zLNOqfn2Du2WQxhghvO
l4HliW4tek7aKFViZOE55eHtAWE5XXKYovnXdKuGn8AmvqTPYsW8x5k8RfWQ3XSgrdCshnjub9mN
0aUS2RtIeAtkYpVeB+YgtXH18967hPPI15+uWWrZXVux/8m/Y8GFhG8fxHmKGF3JtXrUQwIA2PVG
dmH9w5q/6zZ7y1mdOVqIbCno50bTuJqz/kkoGZy2bX9cMsS7nx50e5pUunoGRSU0CrYDXkDMOvHS
EMvXCTrpmcVi5UrI+4Hoitb5hgXYYzpPXarw2Be4as6bVZ9iMzfi/uz8zrzoH9PkRKBhZduwTiQb
61FlLtzJtZWyHikVHi6eZJQjMtJytJMaNp3dw9UApI2nlQMM8D/sfhww3XtBRGtkf47eWmsR6CY4
Olb4QgbL1UrOyB/GWbhY6BO4SFQZSJvr0btOObzsXStMu99PGT4F8F4n8t2CHONg8JTzozEbDLrB
UH3f09+TxMakNumiKeUzAM6ybpIlKlJkoo1G8w/eUSEg/vkkRCKrFnJCEkMoThav5riMOOg1Kj8w
v4g+CG2x1tu3MrdxHhb+pFnLxY7IAMVnX9cFAfmkSuT3xMpdiZ1c3u3lOBjuNNUIPwfGRtC+8ies
ovOK9sABctxwQWRBJc/VCMjRMT42SLSrguoCPQsXxB+qEzdk/tUqtCqsPxKJfCNZbULtDEIycFIQ
LoSRWcUy3+8YEGc2/VtblJjMNzYh+5yQDTHzDVoo+HzGkwnEjay94PHJe+OKg5rgNPdgOFqy3jYY
2BzIZor5TsSV3HWsMXn+1VOw2NWJm4pu3fwy5ICQcFYaGktQYMaR8A1S+N2LEZ2G4YqQWuTUchgf
3Y5Zq4YGUmIMXw25YIhkiElY8N+al+wAjq9MeLRFGajMPosoLSWBhYJKL76VMFqLvgLyBkeJVYRJ
D7puMUbkZvmxge69MSWwGOGsSL6+5Xu3ekSDraaRqmOo9bxaWB7bg52Cz8GRZM/SrOnNTNmwjx+2
SrR2pvkf+s7evxt53cLR7zUFJlUl/5KxDl5TsjpJEwY7jVA7mam+3VrGOc5sGgs0JDYbc8B2dTjV
9o6u7jgRDUKFCxcLNuGKfiEFkTpHeXKsVwqaJJepxHR7EngHYoVrUFUTjcgWZQuLYxpAK2HkMVpS
eFzH3rUCbcJrqICX2Eh+JC4viHXhY9VaLNWFJWJ9Agk0gD1cehyjamkiCnk9idSc4VxYQO8nxoH/
fZ+r/zch6lm+sB7xCYuWoFstHU4rsM4PJ8PWcvw/vhfz6xbdeAx/9x2PFduV8vH1uFMxibJ7XqGL
hH8tO8Dj+/0QYu++CsHKdDj7YDzgVXgOVRr4R4fy3vB/Q00BtaLgz5jv0S/dbNdDIVFYn+AGv3Fw
2m3s9/M6iInxs4e129qo5i04Zpgi5WMI91+VjwOg+RC41qzR3I6xfkXCYqo6p7kZgBoGlQU0i+t+
7hPHf7kRrhfOj3swR2sCpu1VS3DkT1Kuh+rA7IBqnHglS17evd30tMKp7GzWAcleCfX+QhCqKmBl
EPYBotaqIejnd0jcf9F6+TicDbbQiX2yzVpFDuXU3TcsHYrAXgf3+ioDn9DAiX7+8G47QMg3Zg3Z
KmDdDsttC2V1MWZ4oWdMpqfayUC1z1CbM4/LzD3DQdlgSTPp5AUGArmB6Ip9kyHuJTk3S7CCuEmB
GMi233rMA+jqnkN6dOvRDydNUIt/oJgQWby3a+ZS37XvfyqBThxWkPXrq0ziDlELf6HmZ9tct9Fq
//d1Y3j1zOpixIiN7f6iugYmPw6Wq9igCpV4fodRiBCAEmNr/vttsy0CoUjtuIjXIO1jSdSTBhFs
9HllqO5Bc7mNq61sWDhh/roxsHWJDC2ECExQRnFSGxbFyx+WJ6LZ4VHRwa1K6a/VBIi0CwKb0j3/
ru5S8/71MvSETOM74LtDKvF4+QRQCZb8Vf1UxB+/khWS0bqBdNLwCsgKwXEv1imOyPCv6MZY7Izy
8nj3a9/jCc6spsj6hAvGPDW8ugY2LS3fvLjR28P49Vxpp7rSQYh6JMhhPdE4BO7pN96J3m8Y9sFy
8zCHaasHI1zi8Fxm5YxKXz+6cA4TX+0AT72JMFN8/4Xhb35Xs59fmypBsd/8a/jv1wHVFuMckKQW
vp9bLR7/LLj3wWryu4XebowxoxPBcAGReEhIQhIHJOjnoM/OCiUcHBIRkzbpRsQtdM0heKWywRnk
DelnWQIUWsN12JiPwSEtwdEEolYwFh01j5RvXLQiS30L35tuFBmsVzwcVIydp4dt5hiKh4+cYMM1
5C8IcygcDhj2XxVjcWa+hnBOrVkcaliwPZay/tWTH8AYN9CiVZlurTQnUm27Dc7p8za5+QBPWt8P
b3rvH3G/1i90fOqU5s8wzOQro1OH68QOgRBLpfZbzywLSF/odAN9Q2NS6rhyvij2OW5AKFweR0zj
78+hVJGmOLKj/jX5yepj1OVl5OGLpIEn1i3nuPFp0EIPY+Ryj1crhTv8OeZ/YhLX1ijQct1/9fhb
/zlM73tg+ZOUC8Gq2lWvFm2JYUEV9PUax2T3hU8ndJwzJDXQgmU/zx6QJ0PqmDmW5SQ8o65jxtI4
kuviJeF3ggSIcvzZ9bAurHKRROYfMz/OWBf1QgyOcwmWI8N+dILldMpqcAy7dxbHFDZp8/u1vtFv
secIdX8+pJZw4TVKJS3BBJqzavHbBwmFom4R91zvkYg4bJPusMgfJ1ccPT0qK0Ci41hX/OEZTAPh
JDaO64q6sNuwY0ARY+22WcyHwHb5GIR0OTcIuqR8fj0+3g/1mJ3tbb167sJ2Cmrz4TdP6WeJovlf
3b7KSZtXBCSCShUYyQtRDP4wakQWVQvfbU+9L3IxF/fzvqEFcWggNS8RSwk9E47ny2Co4LoP7dcT
iWpwTlULM1Q7PmNkm7AXn4LIItvpuGLXOG905HmG+1Aam5Uribcgi8l/3xBBilymnOgThlaN29tx
oBw5J329tmEA24z/9Grcxj4lrHl76wQxHUhtNZhP7vQunLT3cY1sHJxIpNw+aFcqDO+nu2+dyHng
8AQGBB4koPT0BoMklJwOS0anftR7LyAPoz/b6CepPCp+YfKgpeMDEVJKZcOknnMUifRcSOYIlS8v
dDedoYCQ/c67IDgSaLuCOU4b9yA5/soalx9bcgPnWI5m5tMEzEbJDHNNLeQyvbS0uZVgNUiY8dJY
K/w6gCqQBQd2FrUKQhM1A7yQJkDwm7UkvtwBI8LFHb9ae/rfNI/Xlb2UGOQVNF2xj7fxseA2ZQUD
daCj0gVQk4ox42EeIl3CXZVyCfduz0Pp703MYXoJwMb29dThuDyam7/jL5jiGOvYDT3hjC2+N0Ln
qQM+bZ/Vi40Haighk59anZuSQdHgG2D3XAm8hT68topLLlzdRLnsCkMOY5tUrL4VEBFFVLCkHTDd
w8/+x0d8l38ra+Eyx5IiasYVGKPzx66zGOUtup0M5gZlES8tO2nHII0ME9nGiEOcOf2c31pomKx2
/vv81W7bgvYXxA2bW6DHpPGOZOXgpnmtUQduywgU/J6bxDpDEC6c7uEXH5N/M6KHue5ipwBOsPAr
aQNqmM8MUSDNxGyjwLXuL5wzamTpv8XA/O9MRV49SKT1dusvOaWqOA83npy0aS9w9JJn2rMV9eL+
dSzldzdrvu0waRxpxkpJH9DAAZzIlL8itDHSMDFqxEtsLt4TP+sPk6xOxdNg7CJsCCwT7g1kXm1H
Ps0eK2j/QWhBEypQgY81ORqNRd6Lc/pMLsfazCDsAkbcRGdbXbDwoZhHsHDZ8yDGmjI09FBseaWM
BM9pH3wbaWtrHzl23KhHFuGhuGKPYdf4RnEcLFAp6HRmaUZQVRfpYyBS3dJIEc6fp22LreM8ZApt
Ch/0WLj4c8wKFCgt2retkYG1D6U+Uw9ZUR5rgqyhDIma2pnxW9WVHTl55rn6n2Ey+oa8rI0LpXj3
oan8+ZzsllqPpwfBZd/gB8DT+Vajb856c5SWp1dRoxzm1w11WojLnY+QyL2Qn+KjQ5SQ9illJRb/
7h3xCN74YvzCGsTlqg3WkoU/28lMIMOt90j5s5WEtnPf9rbeUN5n9838OHabweF0Ps4VP+mMgYk6
biGYLSyPTdq82ODwyAShi/4vh0r29Wjbwgz0FXYoQJMHNHBFHqx2npscNLHKJVbxY4jDoPlNYzHP
Z17P1WnZJ9273P1ZclrSx9HQUDnQJphaiHlH79d5rsoqLRZZbMFbtX0lhVb5H0tAOIoc4TkbRyVy
EO7ccVg4dwTd6CmYHaGOeg/ZRAnXxU+2BUctlUkr+SsFa8M/IZIaHSLAwyRXy1o7PNQy/ozwMhA3
16J0nGWO0sDy8QdaSI+7FtPY7CF2nA6K70FY+7ah5zCkfEjOyT6o+GQX+VQnoWoFGARy+0KoOHCN
VkGT0oa+SibdYi9bfX4bgn2Y9rlxXgURH5UA+aLihbiT6iY1ygUd9VkbBXNkA0Qj0YI8+8Ugwjw5
FoHYUyeyq3dHgvJ7doPdxhIPheyUVKHhVdIXJO8Ylowg2Gjl2TcR4z20bxtbf46wqLjYNB4/K3/H
WowjZvaAWthCqkCzcmeiScMxFKGJIunJ6HmZL6ViddV9ZVVHsyWAFsANUFzIU3Z+IbmhaIaKbocu
mtw9AwY81OSu1wVvNEH9UqKouHZfViBp0pjtwfyz+J3EcPT2elVUpzP+mpIHsT8h81QiiiBCRpPs
nrTz1mhoWQOb7IuKlrx4stMdM0ur71cSqde7VMnJETSnqnZi5Ki27vBJzvXKXTlcgfBacQfpUarO
1rKjbaWNFFMBKMLMHy2JWrg5bNCBwm/ALkr84WijvBK8zh8gpPhOh/YI0PeJjw1C2xjNeWrH+X8v
FCljFb7QQ9u/LXSka+hYl5cTn4yUHVVVPlNArNamyMJEwAWSCvOlC2aEmXGbDIS6+WblvniSqijh
HkhGbXscMGNebgwfdKv7Ig9x6p1qUQ5P2Jl5NO1m0aJ+y6udnGiBJXcUHBTI310t3xBeb3XQrCuN
TlngYqGP7SB33f3dr1SfaqrlBBBPf7y1T2ho26LO0BCJVD85SlPQZDn8+A0lqRDt1ZcXWKlBl2zw
LTB7WQq1joodMY4tY/VYshI8tu0aszuFOp5QGjjXjP3DrxKfGz6lME/y2Ovewqre60/Dm1Q1yhZ5
jTsw1mKE9FRuERBsNNCLX1cHzEJh1nhoU16OPBij/ifWpP+Cr2OboRQDLrF/ULspaJoBSUsAJkUp
aaA4YvbELdv6O3ywmKT7ISWBg3G4SMkzZHUI3hRIZIZ/B5sfcK2pwTPkkF/oaDm8+L9ME6piA1U4
0dBZw89XqroRvnl4cbh6RPTooSHGA5ERaiT1SgTNEGtt8hs/AoVOIV8PkaY7Mbb6vfRfNrExUSbO
mFAIjATBU+PNucke32IzCv9eqnAtuJ+naxxKaF+16kS+nUgfD27MvFguHEaUw1mtZKbqhgYV3J9z
QizTAw3Zx0iAk9Uyg0srDTlN/aK0bcz71fMHjrjsP1GySgvaqUzkugk1f2NFdpNTqphFyJW/dDpT
fZTZHQvPeGZBkroQM9c9ejC+8pPW2hBSWSy2ONSKVo4DeCA3RqJAussK1VG1z2ntfBetO8UTa0kT
ttXp0ljORL1HQK3MEhz/DCHfOzK74zsPDryhutpxAHs3K8MOQ2JiTBpMdNDZfsHN+vs+r8dE7Pf8
Kl3FuL4f5yLC9wBbN9l/k2yp4IP6m7l5PGuHv3aab7+RSeOWhXP6gIUyCAh5I0UXQNO182/jCuSM
gORQvKPL9pX8kewbcC1zcgLpCUaf6CoMvTMjpzYIeJe6qSUycrW9DB8Nzf+UTgXhBW1o0rZxB+O7
Z72srVamVSbvoe3EoNjk7t6XPSBxdD7PIBwzUmwVK/bZ/1Ui5lUnOeUg/GV3A6drJbMGbguzqbtp
/Lq8K23YsAqk+TKtgUEL/s0EngFASULDtzQXrzE5SaOhJOMlkzkfSvrdDLKlDiNOJf3kMXT37kDS
IZbc4cJCW8jw5lqeNGKAVebRT9g4PRD+m604BN/Y6HuXeR4xbazlpr4RMyN2H3KEKL2VVYGuZKML
lcglkIZVJp6O9I3R/thXX245eWprkmCQ+e1jOU7XUtgizzAksgZ3wrsl32kHJYPktijZajJGNlF3
eU+0KbrdDznUGx0wgMwkB6Xoku4drtvsD9Mse1SJKZ/X80W29xpJM24KQ880N92DAqfqtyqa4rWv
7hkw+Nb0Le0pQB7x2a2wO9FU3VkREnf/HQqZ1/vfUzG8Ghaq5n3iVL3m69JgLEyBTb/o0oN0cVj+
5yNqcwwiCzqM0I7U2tmxQ2RA9rRPZLLvguroYs2aCu0UPF5duOzVSP+PraEHaFB2NX5xK7/vR9MB
6IqcshyORkBX9f7O6Mp2IVTPdR5p/EFuqnyqDmC/b/1EHCPlE/0Z2wTo/b6GiBfY8tZB9D47yXVe
i4mYqzt1xalb+7HkDobCtgz3yqxY1fe+hW1Bewd+D9NyKoTOK+bKKaNqUJHmLejyF9SxvV2drfc1
8PNJpqIUXOLmRHo3tFLnbcLfnEnf5C08tI0Q69hNtBz7A9+noOc6fKFytp3itP2yl7EUsrxJcTrK
9b+32IuD584YSp6ynRqI1JBs8A6Ma5shOGAFYREvsqvaKkH5dHwhKaELve8CiGZdgPTCE3wo8BJ0
9V/bU6PlKvxTNumxVZdY/YrQFcqSZqoj3kGPSYOMBECLOyc97wTB5Wya9cwLJ50l9aH6St3p3yEY
o3H2om6r33mF5/bdFLSF287JGONmKacIaVAgJpDB+3uchEpQn4ZihvkSgSRjBO2XuMXjt9ORv26/
Yy+ITI9/y5+F8UmblcmPN1/h8YZ/gMESbh1qN9VK+dK3kInKUDd1GPs8cgCrWISWG5Z0t39gpywA
B6ZCLGt/7R8a9kAEZqJsbNpW6GUZ1LLsuz4qIUUxYJOFQUEk5a3CRKz1Kqt0HG/dUF1cfEFljjqF
8gI/5lRIq6MhSAdvhwCRwVaskgPTq9sJoaTnDOsAnX+4hvG0lUqEYZcB9SwfqIAvWaB5YXKVDCXJ
ZQBhk8+zrgrnCFDLuBDcazmsqIIh06U+lyjzs6yrpopuidP5KRRuEWgIRM6Zp7kFv3MTxaTWzFA5
TiFDoxz6ARA+nzzzd9CPz7/L2lsm/2IznwcFltgn22wChGnZmFg+a6szxuCUPyekj0MoyQlrEHQG
0wp6k4oGprwDDToUs2V42I9sCJU8Crnb9xTSc97ne536MpXjvS4X+QLgVdGLsAfmWXvxI1BUORKQ
B8l5qeyr3sw705Xn4kEmmKio0KPdjZHuw8L8wai9OT21gWIv5ij7SHpAWXPnjWzjpgGLUVLTGSMs
FSnAs9bEfIwvNrZ9mcC2B34uK8IRnZtxKwbavTIYvCd01Zmb8jlek4kq+s+OELXosLj7Q7Sc997t
jywrx/SaXy20eU609ozgrf8Dcx+DBhHrTfMQvTTMcYklbiNNizoXGbaEddP1qSBwDZRb2RjJVYrW
UXXeFjoHgx6ohZTQxW89LnxY4xkhsUINgmNZvA/QhYWgSYRy1hMDnHRySWUuv5YW1jHFh+mP/Kfl
vuZ+WGGSEwVDqOrHBsvXhC+FnE5hlfwzibWqPf7U4mGDMKA2zLmWrmq21BzLz/vD8iX0Qj7Nedng
rYcJasJxJ+lmAScjujMoJgAsyZfkixEHd9l4DaMF4SjMD852iFpukE+OX8jzmtF4/nDYT1IMSTWD
4yN+OfCLdb6c2fatGIU8NPJEvDOjggUFeevf2iXKMv6Du+UQvW2FAmYvfSgDLvs4lvMWIPY7k9Ck
h5qrwtsUBJ6BAnkfd1/YrdjMjxqyz77UVt0hOIAt2SB3T8kF1EVnnCaYj6ksd1urXj8ifkn11mxE
5T38G1linwV9r9p5ZOeL9bq91V+Z99zrVjkoZN6zVPxRlj1BwkJxJpAJSrIB4mFz1oyoC8+uKyUV
gHNA+Y64vt5xlN9G7wCay9DuOgHI25s01dM8myGaM86ZdGfLs73IDr0giAtUxq5wYI9Fbq//hfa0
8DMwUdw+GjT4SX19Ud9J5o6sGhAUq8loEpa16CNfLcv1pOPEji48REVrJZ4UssM/aH4RfuV9YDeW
An0jbgonmj2zVstdJBc+gPYSlkHH2yZJoTTTuXVYRN8o1opQY6oESsybyGJ+03Tdg1eDsgWjUvw4
MyvupktUjCJEnMt0G5FrTx2D0pwhab+EMOgTufYw5NJO5vGuLW/te6fkGn0VcOcZNx+36hyh52y1
toNCl8PSGXmh/jdnUTU7YqigxVu5mPmJMKO7s/FhdqHP4SS6PJzsGJxPl3IGrK18sWigNxqzoAvf
rNnaMQSSGxOHLWk+aZxbWY1nbWwasKo4ZnwREalLTcpf8suCMQ3nD6p36jeWNHuKsxfvBg5EcrB4
wuwcg+VbPWLXh1msjyY62dyxJozqjnOM5A5x40B9tv9Ep9MOjxwAIQ6E6LpldXVKjj6Knbk1lMpI
C8Q8qm+j0aeQ+2HiCGxJ2Llyy1l5sFQhMxcdSiwFpTQLUgEvEmXn8mo4Z7dHm02MZ7st9xjbeRLV
eH3lTmJxd/7j2cPCTmOBiTRacASt0NQTrF8GDHZzKDw17QziPqnWeAgKaevn42IUpKWbtobOnuMG
dWQGMl/Qazo3/vpchz7wDkHlc4S3QwECv8mCOvOCOH0Bmzgttk6snVWVeEEro5PkLmywUtMxcsr2
vgh/EMdmwUUKPMI9umcOu/iSvBAQEStWwVzQZVEV0cRW7XpUKgIvJIhtwcz4gv51O3ANfLB5tJAe
UWfOJ7Q3aqfD+xQ7FKU+uvdlfQWdqG0nAbxpj9qNv8fGrdTbwVwJDsSi4UF/SQ0pb6sEqBXNtHYg
aJGhl2oQlhiU1qFrYwSnr9p9f29MSmvOs5dbonPd4CUVFeRK+QE4RvNBM0C76q4S8aOspDOYMFq0
/nUPO15bvrYDU8vB1jsuyAWJ3L2j/OQpN/Bjb1CXyBrRRo5OZ6TE7yvACrB6Qdo3vtoHaQmThkrD
8YSD1kcw2/W8ykoNuGpsZX6strPkxK/wdOcSFEAiJcH9Opv6lgOq9mlSJnSw76bWtB4pjx684pgH
MuTq7Y0je2alwpCwaDQdmnuCs58y5uiXqefqF+WWaLSEXXkgW7Beew7bn5i1waI59Oeso/hkkbln
37iliQD9Y5Jy3jTkRaIKjLvzjyZPO8FBukA2JKDHD0VNlwe10T/DJ/ZxFrL3msZo7k80ttxy1+7v
AhC+eAKTDQfl1bKKPzeYhtpyGCL3yRUX0zxajPz1sxfjaNBlE9+Eo6Ld5C3gNv6VKdzwcHFYSsOo
5nb463ccsqlVMJVBQIgE+QsdvDBKr53E4xGCk2ZOUgZs2b6Tf43Sqzjae7NOXhstn+aQCBImzAEf
an01GgggiSpQ/TNwD0NL+c9etCnwWzqJuBHPMr/ZKRykPA/kWxg70VUT00nGO91osHKcyu4l0OaV
JIgzyWsNNk5Js3+gN9LC0N6KLYh3wKyPK17WXCi6C2XtBlsndAIDilp06fBtcsYHwwn75E8CrLLn
83TB8WbJ+l3eCclFIJCwGi5aawHYYNc5iTJCSfCaDNBF2Mp6kpC8GJh+6rU/icLj4lAIRRsJ6BNL
OLaUa7MuaNE0iy/EDDFozuOQjNx/MLop7g2r6kqJwVLVgtwhMeRtQslQi5se12DHawIC2x5ka+CY
WY7xhcr2g+K/ZVEaPU9md7Z0oDv0Hs1bWEfMsW4NNGzvnRl6utR2T0WdqcvhkfzwPI32oQZ+vq6g
yiBW+exU7g3i4nmbKOt+yBV0D3Q0YxtaLFohBfkMAo+V3IMrj18H+/HeQLovxm4vaNOCDrQ+yhBm
3slZ4HGGfrdqHFiNIpYhhBjso0NdLJ11rIOByOSBFKrvPE0TxSv/meQuOUDGBV+vEUEUq0O8RHEj
YAnNOUwp8CAjfu8ZQpbOtfautQXZ5iUrWiSn/89KZtTG7SRrj+u5Ld6OV29Ka4TN/poFMmDt19Rg
pGPfbixdrF8zpgMc5kk0+2t+vYNp2OjE2neLNQCzImL+ieu+inzBdatLE2n7Us75ubW7hat8BfZB
0W874Ne6wV1dgHhe6NnGIwd/Nw6E+Ov1hEFfem4yOeZziingXQz+BiPNgYWSz0PygqTJNb6h3Uxv
wNft1n+t+iWuxXbnQJ96eyIkyV7u+qze16DLJqcQxEJIBl0HVFUhRnA3Q33ZcpPKJ2aEgOWwijax
7+gdeVpb+BIRMC4JF7r7V/IXsw3PCMqepV3lQQc+KV/2sqNLdlvMhJSFWNDH2QbirpnmyHR79C1g
CPRfa1XmBXaps88ZrtDG9Y5D9G1DfHg0OBiADcfccXRAivU7tVMF0KuQjKJr20Mn8iEpb/aRQAgs
g02vwNz98AqmXkeET2mBO1zopm96yhjZuqcDeV889SpYRGTJpK5Q/2pxdmUefBZvtxwrKKnV23D5
+ZSXFNORR5FCz2DRoGy4xx2JJ7n6HA2o4qAQffl8fdHfXnMjb1W7HSRGg5tUd3n4dnLi4kh1AK1M
Leo+XVac7GWyKGrLr0fMGyccwanBUK9SatrCY9Gf2MTWwRnd5ym76J3sRGlitstsxi1DjWPScPT4
1qeaMDX59G5Ae3FprxaLCoWTHoCDtOXXlCgcH3aezOxD6QaSsA3aZc00VFwfsapbMz3DM4KwXDsG
I0uqcTR/R7s7u8I9O2mI2b7yxnfHq9EgkucYgtF+7t2ShwzLJg8v+HamBxCloL6hlXzVx3toTaJp
lo0CfAGRy6jbWCei1+Xl3rrj6B+pevzilluWU2sjXxG9vMo4BwrI59tbJm3sF7rRqnTNMbxFU7ec
kV1wp8FzIURlHdTY3ohw+86agJDNEu1RNCpbtR/tnq7VqxY99sVeG+c/uVWJSIM8gbUpIlUnDmsv
9f/cOxWtSwRVw3zIPCkdl2ySFDHdN6jvVEBIpU3fX1sfleQeYVigIuVa//H0sCKr2XH6dwry0mYp
TdsZatAQvv/ETAy9XPWSw4Bf0IHpt89yfFu0mFweOqgg5RDiwjVTL5Kngh2/aWAgTcBi1OGxbo7K
rt7Xd0NAqdRYsJ9BAtjGxOF6i+OnbJBmBqGMkUaoEkRSp4X3FwyYLXfsqZxT5bMuC33arVDB0AHT
N2o8hsxfYpK5IAaRnZ5zCFVQLiBW/FH1mZpS5OkF4cIv24NBZtrLzEf/Uao5OMrTYV9OM3qymJtX
WBREHpfFk+PxQKMwzsYeyg25MU0HKXz0uZ2tyu6Ry8EVvwRAXh0WcQviNskeTmJIyoolO2pCb/+b
bvwA6S+ARtmHR3kTc15NfOtsdKjE0r6YKY98IQzuXtOVuJlYr7JhL8LcYBSvj2HajgRf7AwhYp0i
uXgwLetvwrXD0wVj9fiHDe2fEhGHwjiwBa3/FUGCe46nQBT6fJiJTL1EPcyYLE8mx2ba0yXk7XFn
KPST/3m3szmdWOTV0WLEP/KhCe+WW2fie0byuxLcSFBKN2ZbIGfiDtksFmLyn6E+liZQqwmmYr6V
l7qFE5qPHeE5mV98Ek8AINO8w/J925HfgzBBgHw/XquYp6Opz1NfMbok914r4jVaUgzLAEz39lfQ
ImgB0FQY4cwwMTq89IKCA4Ouf521h2YJUO1LfgghhbcxPPJQmSFAZQczUZB36pFzV4DMlMBLYb64
PsFXD6ur0ACZz3qXupBLZI60hsXd6wxk3lkA30dWxTNVpHulbh8gWOi2js75w5CJy/5zrZ3xBUbE
rpfxpN1pIL/TM7ylWkG/VqL5PzVe7IHPFb0hadcypxHCB8SFokPgiFEqsgnSSjzYNkAExSWILr5a
H7soLmYkDzkTl2tURQ3MFWfDl/3OINGTRL21rFElXFM8uYt20a9ldU+J5TeijjXARxKeZA2kLo8T
2d1xWb/2hIQAHnRkgWeMPcndQIYPYSvrIypO13HwvXz3+Wc0xbAUxRP+qnKTepKY8KSrYXHUzems
93h1Mp1Gw1t2ubruA5nN7XvFqz9ckQ19xgggOa/J3QfBlik1RhLxnZUHPduimZP+heMl7KVqqFm5
HfDZYrBKnch0C0p3lKoYdRyAjj756VnbzxV3BokuflM/INU4VuuwHK/bjW/Rb5HEunXaWvArpR7r
k7r73KigbL7yGGTt11tJv2IXW0br7FOXsSfx/HDEk9PL7uBSeJUql6iCIIDIAh+WFN5DWgL7cNeZ
TIYurH5bORqa+csVZf7845yqYhEZaLcyBf9QyPy+A3jHiqPsFFFdDbeBo3LJZNcXdruWDrJ6wiYs
YK1xRXEGua3pYSF4/RGB43L+Eq5tAQSoVrtyXNldRenLfltOjZpTRlmkUZZGyPHCR985F6omhi3p
djJSDdOhArvIuTUMnzGB5xVjlscarhmo2E0h3EOLXshUgAM3gKyOvd4pL6jyL1m7XoB0zqHK98W9
7U3D4ilcyzANJaIMTtppjx5Ba7S/nfiYqrUPZRrljE7UG/k78OhZ6DsseNn8tFml4TnVRY46W05n
emOzCfDOKwDUhegd+auhUgngXL+SseMgtXw/vhJDMUEb1dp/3Ha0KVG6jhsqu91hXtupEEEkAxKE
YgeQdzcyHcCRQNqitqOA5aUMViS/440I7YJCvcRq+M/TuBd47qmNKUJdQeibrhq6eVc7d03OVKvn
/g8owoZN1F+WCXwTuPFw3IB1JYJNVn4j8+QYhH9URnjsH1/PlnjGbrdg5Jk0iG/uLXd3FWE/Y3UA
80go8zzdNjIvLalvqBOQ+RArR3SokeMjDJOp4wyGUVB5J5XWqWffHHwX+GciBPChLiuKnPbJuvWq
e8Fr/JEd1+Tsvkiy5qnD/TmH8APZaQFTxoGHGlEJFMwBz7/RtwUSiQUkxBI1CyAMeqFk6ZCyT817
Tcv4F5q+BfZRTFX6rZkbl3Zdfvx1dlCrMwvYNLYDorqAgok45BjxkzyKtFeSm4j1CXtdXL18cPWB
GmGCmXZC+uo4UvXnHMvbHYF3dI9PRd8moz3wTyA+gB8ObcvPeNvLZZvwpj9R9KR37b8tsoKjc8Ww
PB5hfQH/EqR7l2n+0EaYctY2suKW5uXPgRQNNJg/iWVoft/KffNvIhwWDe7KhJCovnVtR+JS0BM5
7VeJywDgxuObAV+mN8pMR+N3z5reTeLm1JAxd5BsT/Hlo8l10QjLVwaVLKak9NbaU9Wx/S4SSg1S
Y2136vHp7fRiHSduBPS2Vx0RICLEATWZ8jCm3S6TRggNkVe43BGAYT3lzLQJcHz+4MdgMAn+w+cm
79eyvrn4dkyfmqKtVZmUTO/xERfrCBfUCzmnZrK7dRq3cD1m+X1kbCF2UDL4AmN6G4AlNO4mDJGn
hGI9sb1nW8QJuRfAcd7uCLLGtVvZvcaO7MLrq4wQsyPgS8b2StQuIdg+kc08wiEO9PNSBbr4iTb0
MplhIZrR4Pv7P3DnZUoBwg8TP6mLGIHy7nUwkj4KjDVVMvqi6T3I+mcZnrkooYe2uGkBZRCicZPg
Y0qR7etlKVhk0F3GMmIIlY2C7fscUYe29KCYj5tuUEu53KKv/ZnE5BMwDHXaEkTo0Ri3Pal3TRnq
lxmHEpbQjUcDhuo5EZN8MrCUAeAcqffbhQZDPLGOx/IFHN7f5qvROeJ06JiiyqbnsEROZP8Ipbfd
THlgVRY8yvVjXVXC71yKwOJOFxy3UZZ1z9HfISu9z+iShXTPvOjAi31xkWaV8sWViG65U7yS1JXP
c6nqRhUS3qciiC4xr9dKPIFc9Z8LlctQvJDXJZfs1+NsNiQZtJxmGxesqvAKIKlKmzKZc1PLIVvS
v4ny8chab9LNM6XXeHQxDk6mvmT5XWGYnwYhq+tGm4zhu8Cdf6gmpEClaQFwWwqmOoWxfvCoGKo1
NAG2kdvQB2CbNSlxCNX71xteV7LXUW/d74yipOYPenYgjzFex4y88Oczd/7R/dppjHk7QAi3xcAZ
blqF29GvuV/8ZTIHIOGzFB/ycNqzAIjpldnB60ibo2AtjQlC7E+OoBSJwf/ykFAVgST+SK7vUuAe
dAO+r6sUV7oqL9DLg8swuWqkw6VpBjx9QJOcs7Uca79XQdr6PpYeegbJ7vzHOZYRz2ClAjF2a67R
oBcrUweSa/2oeqZLeNfDWLVSTnfzjOKh52tJm+1ruens9Tlotrg3YdERK13sQ/r4JUIpFhDs9sJk
lsO9hXq78gQMDgj+l0IfJG67VscesDYJH9hUEGLHBz3vn4us6/mTz8ycHWu1YgsvoTmwB1wdIEkV
4aqwtqo8nvPlzB+n/2/5tmoGLxz1zk+ytdcInmXDSJmOk8pc2WoT1ReqOVEJLv3WTOPRf5VgZ+yB
tVv0J5GfNZQZ0uPuvpOsi3Km0YjVXanOAuuPBxCHmS888v5EXcxnsy5aEE+g7DMDs2vH6D5fac+C
xvMWqQfpK35gNNZ5GvCZvsM/BEAWguGuC+cL2ryc1juZqPKmtzWdbV7PKVeQJXyORsufRJxLArpu
F38n2EcggpSFiwtLb+5dm5nf87VwO/P63rcSM5THKuiVfs08EQq9UpORwcUCW/ZgIo/LapzKxW4/
qs0w2HSZtDmVGD3AO2DJSmnVFhoZtGumgmodvQOEjHIgHna0jV7aiUuiA9nM0XZobERe2kT03GMa
AtNmSnW34aHYhIV9B7C7KXAmS5GhK5rX+YmxBmJl4wfTzN2Qi51PjbtIDeNDeYATMvaRxm7b2Nny
6i5s1lujaQwlOdAcQw+nF5yVWoyOUZgcha2vb4rjPIctUXwRhimz0Nn7e9I5lS4nBQZoklRKq7dX
AhsgAG9u08FtI7PslpaqWjTD562s1fIHK+f8LWsMi55/HCk1qTj8jDYbwd2ooED/O4T08gYTq004
iDhKhUGm81sQZpRwns1R4Jn0NX+BCT0ZXiM+00Y2AppRMHTSL6blvKiocRxQyK2hF0FidSrQ9tVM
42uLO+VDkhYFZyE+xoiPwnV8QLtzJaK8yePC7ZZOCH0ZdsmiLLU7191RKFuFrfarhwZgrAfItDB7
wE+Z0Sk3SjztWeWva6bdiFNXVyyPDCB/UA9ZHo+IdnIV3s+63qvCS1fjv26K1hmI85QVCyxyrW6c
IhiX9A2So+bN1Kv+7yrKaKBN2aCZ2t1KDzy5kKFld/xwfCvGlBf+lze7BaYsiVFgcrA687b5VfDS
atwVtrW7K1kCdKnx2W9ruhZAi9oZLSlTc9RKJCXj7JTyZuLPtbX5PQnTzwOgQbpRSjoQQwy7T89i
ZjqMwPcbjJtHYcvNMXPUKVvqd0ACc2JVKLmNsDgbErbFEnpVkb8b5VgLuJbUB7XgMCkODfd3VhLR
/xy458FDQqvkaTuAEP1D98z/wmwljFS6Viz709UqV96NgJrlX3sK3nOORPXLFSYqI1UPhmb2wSQ8
GT6M7hns5u15aClsCurOIhxTr8gD/dpuRuPJMor6xSHFDx0Y9C2w/4CV9ByCPQnuCifLDLUZA6Lj
Gmk7ODcWTkbqetRhyYtD94fuxGaDq/YDv8Agq53HiYT97diqxv9NuR/3mRaj6v6BDjANhbiE+PkI
XLFuxgz22KdxwjmXdeKwmY6qny5KVOU6505ZNYKQUBBukzJVNYrTy+98vs3GGIHwEcNhvSVWs+0w
WALtaIoMRQ5uE/uvu5cXPWZLT01eQPB1MeR/xYUd0DQ0adZiXjIWERO7FqpaqhLW7CacjOxuM9VG
O/3HG66QuZd18+NSO6lUa/GbDMSMU+TIHPQe04KhJcqmvMgONZkjLJGITiWYCTX68mXCtYLVfzSi
NXipaq4weAngna8Okt810UkQU6uQh+DvGgxf8kMvPeHeH4URjzc/1Iph6YInby1Z7JwhNXGbAtaZ
5VUEOYsHr1kNpGAXsdCRbAddMIE74RJ1ipg6tHh2G9sRn9pVTn5tmqs68AxFTr6uuEyQVKUKvhmH
PNUhVc0QzR/qPDjnrKGJbYkV2vqoqG52uSdtbNwJHTQVKJfKzxKlmGInW3vjVhv8dyjByyXXyTow
1sZ/XoFDGgaJdzZpb2RXunp6NczwmqyZjHr0+ALkslrEdkEUrv2UoJPZReOh892IZXOyayEqbLb8
uspjGvJj2ODsnkzpZfE0Jckt0MtPobRih1icy2q852VTVjRvQP9Xalj/9oATJblG3T/7cB1yrADT
Ng8NZs4SMFMZ6FI6FwW8XNXOmozC7DO3w+4wpOP4sZ3WX5zUb8CCkGcRaGFroMdcoCh6ZLN7QmEu
3rREsUHQKHFHTwmlT099c18XCDdW53KEcbolOPdhxCenkHt+3aL4R0b0iTkttBpG30pq1pw6o7bx
+ck7ErhkdC86my2U4wdNxHTfGWjPyyBlMxD5sEO8LnTUxzse9ArehEZ1KkzzL7Kw0s6ICC8TykZ/
4ddy+VJuJhwFNgkKh1j6klu1NgUBVhA/ym3mdGXO/YBT7bBVhpyHZvXGqRFuNANJKqL56yuedrV3
ktff2bCyJII5ZoHelLOP9nTRL3UjiF3NxrTyPg/x+mSWVQ6q/pi/mGSzPbmvToT0NEEJVy6IsvHx
4R94dceqDoMjWEIvd2tbFtgxCXnfY6MdxZDI1wHm6/d3mMliktsre9aaWatteVCi9ozFv52huTwh
kZMwfMuFmFM2c76Cp2CDe7FkuC2r7YG7DJ9K/hpWdwLR39ajnQLb9NvaxzINBa5s2TblbLjrhdLZ
0/HnjuYIz0tU/8lyONO5i+uixJdk86yepTY1TQJz8d2LShd3EuVnKEAtN23nvPw2NR7oNTUJSqkk
wf0okB46V0ewMAfau7uj7BVq1evic5Qx7P3Lruov2ac6i8vJaZ10ot0c/ZIuJETSxu/XPzEthi6S
FGajOpd2lQd7CQml8MuSW0NyWe6i2e9yYGyvz7Rwu9n2uuiJYVs4axfRfy10BuQ6c5+Nzb4LCiso
iNpg5fyyoqHV7WcMtVqClELre8h3XdJkp7wv37Tv68C0ItS9CrqDcK9pp9tvrSAGpOSotTm5Xd7s
u/uhn7SoNloQS2YqIzbGCfL0m3eGNjHjl9n0yH8lJiyI9veGrxm8ri567C0Ad0BEw4eBMqu4PsRb
bCd2AQv0T8lgdocCxreZ9J8K+XkFzWA3NpKPcjupUcj1bDeub8CUWzmb0BWdsF2pKrVWmBMApMCx
y6vQpdBBdLg9leaqhm2jPuhslP3tercEYeebznHfloqY1dxeOvnGNKFl0iT1at/Upbd03vA/yEAv
3iYgA3U9jo26abUsuscFZmGAB96zOrL9BJwb4GUl1WUq7qh94QW+H32mee5DHMZy3e//vhYvpjnV
71D0HtrQNVdlA7R6v5RhkpsmFygCf7b8DZnMQczLt14F7M0n87qBbAp/iH5t0EObvW0Q4lehoJVs
vQK/sqFwD45+g67BmW1y8fJBP9+CT0MW0NdTSD17cWb8eDuArkpRcFa5gC3NEGC/BRvWswjU9QrB
H1gPGl2IehhgkOpZlkwTGCLK3s9cv0EO5CeX1giy2xVU+VmG3X1iPbkg8BcdYRC114IgV6Q/IALN
kwYoz8VFB1/z5NBA3JL5EWYIKu7xZSSdrnrtS5DAt3DrmfPfZeu+uzjuedOMU3WadSiFbzcOaHIR
fJNy0QnjNzAUZKRWxzuefh9yJ53s2zQW/8lmZ8lFxIa/NxkFE01D81dUiPg9muwxHTtYe6eTNwYu
WI4HiwoezmpFt/8FTthS8mU/zwppDj/n1wwqHDlR3BiUyAfuBgRLYlaxTL5ui1oFBVVD0kn44NqV
BekV5xHDVQbtcSSHI73kqcodKubJ5v790YBi5f4G8vE9KMig8+0if5DDHqRwPtVWdguvyIRUJtrz
dUyGc32qeEq2dgGbGgdzGU0n8I7e03XumC85Pz/bnZyDo54ldNzn0RxOcRVPPB8MSI8JcRKcmob1
ccLsNsXY2NNrLw4tVTmPpnxLBlPeG/LTvFcmTc0j9d1ZmfhRQxahBkoybP0BNtG7W9lnKU3XYngB
LkNjgDPO+esNplc/HDZYfTknKMn1SWmFFrXwW147MscAjpXjpy5Acf+PMAiNdauCJSOiQw8sDlnN
0YCSsowxAV7XK5omkZuNj4ZrnWC9P2WVK7oPNX3wcQc+inf019/b24qeTewMNtRPc/c5FXUdkfKf
IWVt/6lV93jTpCz3uKuzRUb8mE7KVIMio2Xl5gzIOg9SFBYiKvxh7+FUYSxNRkUtENBKAYLEiUTr
W3PRS39Thi6KQq1gUtHRYsXkBS63u0xHQsPTzOXyMs6qluYjvNFi8dOgOjUylPsNhSQdn8bR1a+u
FpKJaSeva08wOjW5fnQgjrJ3jOHk3+wcxaP8KyZj2e+WaYOVjtp30z1go0Cp3AjZTbn1dX0pc8Wb
97jVRKox2MKgKzz9cejijsoXb4hlJ8xVgiX/V33EXVkREMs1Ong3WQtxUE7bkCfLxLnaI0aIwhpz
vzdSzmGi3z6rWmszQ7ku0ZWRIX1O3k9TTCpESUOyEQRcrtv9QcXtBJXLYmGrpqFOweczEIURqrS7
/LY727ygU2+Izf8HVefk55xwBZ4fRDiszYM/obQ4Kk0u+Z8IFyCC09qDw7Ma6vBtUvU4Sj/ioAzk
VcGnLi6vmBGwBRUOQn6o0OlyY6QRHzs1frcBnfFXmPc9nTp7SyOcJXfZT1XanQ9Tux0sR4QhNShb
wC/bTFGpkR7UHa287gZwxiPDJSCUgpoL3YOA7upHSbn4wdQddIW/NpZNOrtzfEOYmRh6VGis16p+
I9C67A6CWxAzBrNlMFSuitxWW6oNQxNvFTmUHZ/6zrMtLkUoNQjanatgEb295AObX280eZDZzjpM
Ifpgadwk3OHBBeqRY6LpoGMocGSEzm8UCUX+XvdPqF50C0KWAsybipu9RHybwr8oE+FUDKtl6ui5
0VG3AUdZ7UTc6M+WeTlHmpLYwPyaPCU1BXcvgUYiy3JDjRzjHgS9rKy5HPBQ2zvM/9HjIUHexKA0
SmiENstBARc7feKpDCPVCUf+ycbjOcsfTr5d/5FH1XDWsCirEv5CSbFfDiHU8cZ41vNeue50r4RO
1pUIyQ0x7brMUhjXcbPd8J2EoPavxYI6dMWuKpGZ96r+sDepQpC+adrHPwjPy2ih2s/yLHdh4zI8
C4YrN7F5b2O0uAP4Ax1MLSoCfbJGLGAM0IspQDqTEpQhoAP7B8AyHv2rrR/8BrfMxNB5BPblg5IF
m43J0afeR0lo/9mRpn0V6LpYahn2Bn+93KpHelwBuSAiDF+DCHWJW0LgTeXvIZc6PjL7roxNZZCb
mXpYCQFWszyhBcZeL5dL6kSFmhS2LIRpoNv8/pHtif5aolCy061VQke4nL5cGxmtpu24e8htGBRi
rjuMd7z5DWnuSWl3n+PUcKDKiwRUTPIfHyXwY/lcBuvad2oobsnlb9ZEi+Tf6X+lZRADykTxH3ZQ
GyzMFHst3mJNoJa8+C6lFhHEzze1VgYtLH54b/RIL+N7oIm1MPfT8iSlUeY5UE+n8x41/aPJHgDU
Gntfpozn03nun0N5ff0QFQnpEdpAFEnhEw/BE24afrYK+eY2eBa4uTuWWj7rUy4rrGvAPOJQeWNY
Fn1DlwL+Xp/sDSTUoVBTDZtWBe3GwSDc+2nPH7Cm/qqoX7Ryl4daRGYy1Q3JMjvS858uC4F/QelK
0YbfiRwgjnH1hwwaBeI9indAhtqs/zTVOJjQ6goOn6+UGZIKiBZAFyEqL0Z0JgMcMNMo0pVK10AS
Gmun+qr2/192XaYCLV+NTHKNMAKpgj/QK/MPghztcw/aySadRrXLdRSYT6YI5ucf66t3TYRO+kO8
1py9sGEcoh3RVX3he99LyFg/6+XYb682ZmzwFbNIeC2a7zGJvD3XlxvZwrwd+9voUc16qiAdiqjS
TFmuuip4hcvqRHa+425Mmk4A9VvAOyy51uhHFbOqaPRHUudQj+2DmvWxOAv7VYmnRoBBj89ygM92
DFaAtpESeApF9VdFEjlatM/6lVeuukmH11FXw1MgDDWuHX6mAtGHLPJrBRedozssbWobr6kCLauM
GYjB53K1im+MxtMC6FEaOGFmxAWg89U9mJ40J6+y+99inJREfsrZxyIHDyY3AXYCiChTgJ3Md849
BdqalCOIlKjQw5baZ99HaKnE8O2FsYrO/nighuHkicYA2KqAta45LRdM6IMVJmRRrSeMLy/TwtpL
25ZfsoL/jSxu3TD8J0Z0MEZN3hc7BM11W3uQmHcL7uW/4TmCVeCzEJOTzmJB4uPCGu58/JuW8L+c
bCAJtaRRJkRoTRooMsxfSkJ3+VCbnee44i4AWX7l+MLa055wtBqyB1YlIZViyfmD0Ul0REH/VpSF
CXYOQXpE7lrLQ/bHwhtPdFlPDG2/ShD3LTPvXvwEOAO2qmb1JWouGtSlCVt88KYuhyzVcuJgX8sD
Ew8UteLUxVhnkw/wpja2J2fvjkGHSAA9TZsrSx/tHITeTX7qrPKnsG6bBBP9q8RLAA/DsYGnzIU/
uK14Cj5unDDMzOI2rp1nJC/Chy9QaznhJSvP9+pnDFHUz9JwdmFh0CV0VbTeCuKY7y/Z8FOEpCBN
NTZppKQnA06Dl3Kf9CTK2h/LhgUid2yX2s/VlYaWPExg1VC5Gk0uQ0Pj3S6EBtZix/Y5imxMdQv1
ND6V83nxHAq9rKEAKKs4HaQVkePgsI1iv3fUVj/LJI0O2CRvdA17o3aN4h3y6ZkXXsVc8sOVFltu
J0qd1R+1bUUJGGgkaa3tBnaCVwRcrjwcsiiBt596sXODROxEGLoirOBZ6t/54e2UuyliJrikZFl3
kxVepYLVNxeJ1Blj+f9/Px612ZpMhICCRsjBGjynFfEnNNwQHqRjRPqTf8lHvh1kr3rxU4PvCOP9
K3WcDPkxtPICbQjZWNWwESoKmoM89H/A2PWPcgWH7AnTsIcT041cs9U332WcxZdaXjJMucW8y+FG
D/1F9xD2s5Fv6KK1UdiOAIwsUDDIdtershWopmEayAW6Hqo7/K8BPu5ietTAaB2rqyhRyMXyUSOy
c2JZbpXEx62ttoqh88uLKkt4PunQa9j/GmO7Uu10H6autK78cQRQnOGS06r2dvFsNgRmvfEbiqan
ojTUMwmg7d8A8UcpLLUbmT7BhXLv2qZPwYaopLdaoBQHCBpzSFSW5GWqvNIE2et6H++zTrR2hL2N
kInLrHw9h/ECBe0CdpGKtYYebFrLSdVfSmxNPg6isXQopiARM0iqls5GzwH1gZTo05R4+cVrREHF
OeisDXdPoNWEQ0PlDuLpH25Br0SENvg3f9Tc1ENytwXzAfTm1y5J4wYRD8v2k7KtvSfVvvSlT68P
A3D0NvwBNt5gE+sNko5peB+2t632+La08FnKcZs3zCkjeerH947qNJYwFYQNU+mgiQvNWtKdqGa6
JbCoWcIn7m0r9J7aqmwGfkyAj10G1M3FN3RGdmlS/DJVflAy6AGAvkznv1QLKNSHau1CIkk/JYHZ
BeT/U3g/UdVQ+D/c41NUHfmi0WMmwuuq06DsXLMDh60nsjo5uvV1xkdNs6F1tIJW2uNlVH42j2Ia
tol5xsRgnKRjCQVUPvw8wbfeNx1NGFvCsBcNNaUjHaIUEpUOSrfOOisejWRDFkrW9BpqV4wzNeP1
/x3phLry2VbnaTidqOSHJup0X23lyGLyT54Z3RpBvIpjEyluCRImuYsIC+7m0sPuFvUZQK6V77Gk
vRs6+B9dfzNDn2STQv9eqI8U+5rm7z6Ipy4WlGkIgZT82EDbUs3AO9xoxAs82ZKgqYiKaS97+BVk
UnLjDuNCuqc0cWiw8Y9c3hVEcKVNok7E0bAwELRND0Hk0GYr8aRQfsePSsmKN9G82SBY8iE3LHR3
+Fry+P9AGX7uGBWpirnZqdV8y7x4n/fA5KXCpY8Mm68HICDhazlcYnznO3bmPDcW5xCoVOvKHAkt
u9gEskI3bBPURMLKD8stonHjpGBSy8x7zOrzCoiyrnZwZiaflYVR7hSoJd9LB/szD8t7zIqDxAgX
0+FhSoNrtWn2YnKcBuEcNcs4Mr0Vw+PnvnbMnnlv30nk/IR5QDLAGrh1jbtU5GZzvDt15+GcAi87
IVKJxsjt7DUSKLpInteZscuH2hoaYSfE86kzBDcT4XdyNZFXqRnUw9kSbh8tohoKHvYmgcg1i+i/
ogO1OoboU83ywKxi3DXhF12wdFzhEV0eeyouBEIhKgDIGLjYg2P9Fn0dU4mv1wtPX1MVmXrsvv4f
q6jagBwYFFU97Iuf6GUF+hkpT8kkPQnh6ZZ3Whf5CUoYqYhhc2TB4Iq6DqpWLd1x75VseiSlsUS3
rkF4BmT4ne6Yh8eyTKKv52+q3O1c2RL+kybR1apDSQ+9qwExaCixUr0ui/BlGrSx1+GrQ1R6mdTW
AB7WUgKrWR2d86ITATO3Nk19oBFtWpciEkMlZG14kqdJiD+ZCVxZyNONcCgP9y8I/xPxz+Y/Og4a
lCV90oPNW5f9tf8TfaLfbQj38ar7UG9Ul0hV6W8RWrZHNLQfIagzRD4jO7SUb7DndqjOS1gGAXYl
4KG+ql4//9ZMCrEGyojLyHX6DZgYrNlMKeJmEQ5r/W/bkhy2XsI9E9Sx+TLcVNtCiod2p7sD23br
7m5l7u1vxrmbJbaqiC+6EIUJg1E60glhSsD6+SUoc2gYt3qcYu2WmUVod7glpebF5BfE8+1psGti
kSJOGfjFvfcsLEKE1KiQK4vgEftzBTnDWGW74zCom+q51PkQFSFD987CMEeXluSyXYihBP3pcdEA
uwAC+6t6OMS3PZmUH3Vn6y2cPnfiXl7ev0/i5FzMFpojv9EPcmZbAtQivnSsHa8zORy8W+qk0KWP
b5nu0bD3mTXv/y6t8+81I7CMGDel1Smlfy8Gyqf63fJidPJLVKq+jn0vZyp/DvXZ+UcHj+DmcCfF
mynLiWR445BpBcOWFmj8I3mRMj1pBWrl4mwle3f41i0cH+kHtjIt4C1YfW1zlIZHYBfnkPXBhYpR
l7Z9gJIck6kprpuP0l69PZDYfkSp32Ft8rVYGF7gr2mAKoOflyPPQ2/9BrSVfXB8dnIdsk+IABY+
Bq/rdHxKL8x/rrz3epuDBHm+efBFs+1AtDc400WuW4inbvNcdf80HEnuVqUG3sZADxVbSqUH4jns
sVLM7zG9tPAOstnONCJOvdRdbdu/pvy4GDBQes+/RrLglPzrv+ZTsGpMkyU5Z8WkC1o2jhMqjX0j
khiPNzF3FNNRqw1VFmtwovBjkeWfx3LeqwklHy9eQmdC4DjonDvTFt8XiG7dcGF4HExCw7/HYhsp
IBac7HDQbXsuMJm1EhdyPTySsm4rYkUlzTh//t5Npn+NM0sc9wG5G01fZewYkyqkOHsJafFDn2xf
TqkS4iKvXzpXaXPWyOjIUcPtyVwkOSSHYU+sigzDR24v0+e32/f6H3+UqjmUeOqpZt1HF6Sw/etp
jnm+el3qkm5RWNb1SmYCiosqhXw73r6g03VkJvBILjzI8TxWCD/JGDtY4maUuVFxkcnlGpazf4RE
x2mjTmpt0ExQtkgsXfBrekVF3APsCCLY45/3QF63xcHdE1z1qXatJobPR1cE6HAj/1OX8oo7iJgI
0HdNlSHBaLJsIPAn0PIIN/oyr4ZTi6XlVvUXUO4z2wwyuUjTLP+OLcMEHe0mfu4DoCC8p+JF8BiY
6S5EYuLsTsWreaDsYt4GLIb2mRYtYowQ7U+gn3gC/eq1hC9L9WgZ+kE/Bds46Qw7rei/wzuVqyob
4J/8BXd2pcY9z/qCv09WAZOe5U2GOT0G7BDVL+hBb93ZgjdE0JqinYRakjvVPGLzflKeps1bCQGq
9i4C7/3dg8gfndExcYlH5INPN8czc9KMvIG5umAukLdmjZmi7rh/TLtXEpYo7OS1QBGvls5WmGKy
Z+MTE2gP7mCUCE0eFhB+YisKu3QiBXJo/2Nc/TjTaIsevC66flyZxBqcXysCX8urNoy5zSLGYJKw
hbfiS1L9Mj4cVJSMfpOf5qarSrgVHEOoW3TMe/aHzhq4Lr943pSol3GP0avw8sl+5uZZJ46XfiRA
WTHIEU3TnEfZm89NnfW6qET6SKG5wofQ3+ojXMptxntKcLOJ1w2Dmm18e1pMnI/Mw46NZ2d7E4l3
OaRD0Cu1iQMKYQPC7n+psAdKqAJSphmoX4xfzZorl7Nz5rc29Fy7IX+DU/Sga+YYdbw/tV8zN5DG
CW0K80eguIJ57NfMEx3/97rTG6qEn0Bs7grlpkxzF5RigchY1nQPyVlJZJl5FlO/9W9SGnAnZpho
iCN4sgm3bU54vagqzN0Ho5olYQbk6AJwUgkVKjXuGwC1W8OmDaYklRYi9IZKQpZCBIuHlJDrJcA1
OZcajesQMXDubxXozTSrnbNfWnaPQC+6F7lUXBGBIHoETzwKc9fgNQXUe8ZALgJNV4N5FlK/x5ld
sAFVu8lZE9ebM0Tph+GKNHSJ7Xd9uDKUkI8dpwuArYS+xAxsGBgMkvmr6o+/XFKmz0WAK5+EYXFH
qR53+l3JKhfK7Z9oasHFI8GLpnXl6pzIAq8FcFSsSpnamHUz1z1PVQYTVZiYOx1fkNefxt95i4CE
+1t7XU9MIu5EeQp3ykAz+xzFTvJImsdZyQW5vIQgFFf+i2CoF/9GEcpNOe/Jplfwp2F6xLzxKsje
MU0USQbvckjGU1LaznnjV8DqIAD+c/7HSGzXAD7fe/sB3VryvO2deAgZOeVGv+fzMaFCgAS0peOZ
3bdea3ZxZTWmGG+0kuNag4rsWoxba+Esk+AfM4ausDB8ICiBFiSWbwsiYYQavwgKxFOdmuIvpCYu
fpvCxVqdwhH6MryErCpyq3EvCnRUTCJbCSjqsYyJ9lv134MXcsHlbmHLJv3BUaWRZnLpJbVpXLFW
zCCq3WpT3jqoTYftHF8/VIwEgd1wbpuCoA3RRpFJcKa5J+SeimnQkvDQ4jEfNHrmA2CJjsgecxK7
m9BWnj/qUsc8aXOXLRMm472AmbGwusOn+ORbZQjHxP7+wi3QjPU0TmGw3bvxHSL7cG/upoLGCPNY
uBk/NNmCS+ApQ4Qbhs5WvnlVgyY2VGM1WiJUtmT6V25bgHKf9wdF7uXf+jAqgcz2FR+NgW3uygUF
2dmKJ3y9oy4U4gs73IWkKlvZ8Z7EeRO0QuJuUCojAa34X9DbVhDTzgrgJcXkJaR7HSxNnYcZCLcc
DkwBl4SLIKZoIRcPZSmr5crYhRQf5N/uzTG+/9Eyhf4kDkZQN5rJY/honGgJ80bKK7StTTafQcKe
Qa7RJInZHrLO8X6st2/jzs5nwFMfIVTKxRrstGDAVFk+R/+K9sPCmZC4AxM1ivUIUal1Ekt2sRU7
DoDjfPmekSNS+mjBjzs73Ci5ahNBr70V4Ovf7BbOEAjQZI0a8Bs3eBDIAiiTjTxp2SfDDkL+fVYc
40ESONSoARW/BkachqNhk0aU2vJeOHj9foL1f/sZRZ3SglAGNZe18koAFP7RXtQb2gD845h1VSJE
/nflZZC3lFay+uXtc3ww8daL//6radIKjJ+XQ19ZkcyzQkM1eekO9bHgIZgyF407BUfizJ+0B1AJ
UNhECKIEVWXHgNq+LpV5fWqmt+oZ8ZSPycHb5bRaR8XEckpX8CJSLlbPtprLWh2ae1cAOBqhbT8M
StJ5Ehg7P0zF36nR6SMDYrmEOQYDe8ocQIhXyEYtOS9xtT2Ya3Npi9VN9WL1ZmeeB3KqXkTwdlMg
h12W8QcbZNMOJTBUKcAaB8wrWNR22CvaHZmj6Rwf3rw/wOcID57hWH66JwDxwF3JDyrgvoHafF0m
nWTuWhILq0yYqEbbZ+V5wZDNzfTvxy/sqGf3grBBow5KbUiMiPYpwanSDnPvMQQ+IaMUj+iVY27m
rLWtq4sQgGSeb6RWeV4ly7JXwvifR51zU1VpUYyyrTQkyWGGK7wRJZEWOfJ/O9OtRWGhBymLhxMb
NyhaAGDsW2UkcR6eMgQXNMma3S2LvruCGH9UQm3rhPnhPEK6vTFRoz0SbHACcncwg0QdmspThVRq
GdpMRv5hyb+DMcLONouQQ30oPqSxDvjKLdQDQYCCYMemaxbMh4CcJOPn+3QgCqFOQLs69IAxQxh6
yga8f9RgAD4lcQ6Xak9zsk3buNsWX7f4jX4Gzcb1wwqUIRRjIvGgE4qLkW/Lp/pGH8iiQahzdKWw
cbZQzmiaf+76j1b/0OnFkU1Au6+hOLjUpK+wPKxwvV1min6v4kOZGYpRISgpF6wK7QHEbj7ZTdQO
ijQh9WizxkLgHLrGdwVdVNebk0FGg2iwSvEzNHB0yjDVlr6ukDEBJsHI0hnnJ51S7PbozuIiPjKV
lT1BG0UhAdFP59aj3+egL1otd5MXxjb9ernAUFxb78CvXk6ZfZmtVhy1UeKkRsA1bMJR2kKv4FX8
saQ15PHiuqiQthbFgFMoID4HZbagw3ngYm812TYFXkqS93x18xkKYprGe5QlabR8d3s1s4z6Pp/C
A/CsHLpD0Rbr86ft0jgaNS0MXPEeKAuz9Gf8jCp8yY1bsgQKu0xMP6gre3M9K9dZoQePsW9v8Uac
p4wuTcq6kFtmPnDBd8LML6+2q/PDhLxrYkcsfZ53Sk7KapV9JS+/YIJrIFxRw1tVlUnpPZ28+mNz
pTCzdBtq3Mnb+K7BlkC4Jdy3Cep3Fz2goth4d5c1lgDSvoeI2EvpSdPd83YdzY72ZVbgnAEJiXvC
rMri9akRDRW4rcuPK0fNUduydWJ3gH1H6oiH1b0JPKTo6d2D10dradrpfm3y4jlMprCa5rBD0pf4
MX2wF2pSkZbVnKhjthnTRwgETZRbqdwYA+JAkZltCByyJc44NUn0f2D2UwA9kVNt4G0CUE3YjSzy
P0zpIJPExjkKaQcJIhgkYRY0va/m8/8Z+2glr0/wY8Gqsq7L08SnxXQ9/R0aTSa9oaaabf6x5w5b
yVw8fNxtnuMI0JmhvSqowUiosxY3aFxNpeiOVQdv+NIv+9u8LnDsqeZmpGUz0BTAeu3nhgOgyFFk
5b5hAIHza8pmjbWZfJt9AiXMEy5iu6vGm7ke9GApMiI1AX3CGtTIsCPmh7vfFsZdwi6nEdqm4QlX
dzXV6RHVQZ3XFFluiqeNwRsYjOeTjcw9NZ142QSWtWbfjhwSd7KEyi2M7jEpG4K9Klbj/31nBsO+
wkz+CgkbbUCrEjFWxlV9YKFXgjImHrAEeZCnX5Xrilx2U12tJ7nsjzH0NIMqLxfchqjP92uhyUwi
zK4A8lLV1PyGxUNu0EfTvQF9+3bjJqSLkn0MFJdzHgYugFbZlBo6L8loznwUM1X4FytRbDrFhMs4
Sx3FrbOMF1WHGBi3WHoaC/oDvNXxmkWroYGotYo7Rl/zkWxm8sinLN8JyHycH98GqWVJ7Zvy5++1
RGY23R6b+iWb6qK8ZtieBjHuy53m76GZt2X9mcINvz1laXQVAIWxxr9FxEuPwSKNkaQG9k2gzn9r
cNxJVKqQtblcZzyQk2EJBauWzeqpaQt1W+P4yJJ8UdalJL1rvuBSMj6w0YPmvzii9JBKfooIB0o/
KRrxdmrZwUHhQQSUXjJ/y9MNmcQeEw9YN1ztZeUFcEZep5FFrlB6TUcOZuwtzu5MAHPBrfc6yBo3
RLHuSzF1RAgGgV4cxjG65mB9aTWR/fV3vphfKUM2bs/qW8h12LlNLzLVBjifKrdtUCcUT4A4Iv4c
wR3Uwto6TpoMJIHgqsquXTcj9zWXeihpPoeeiRvwVvx0YxN59d/1kVmhULNtfnOvlbWYk9WFVs0f
tx+ea6tJDF0WB9X+R2DXyxAvY/YEIalM5AoZ2h+yAIIQJEeUeD+dd3cq6NAMh9v0oU1VkDtGd7vX
VYwDIUaIuexCvVysfN9WaQd60x/0UW1NXSEF5IOVfuwKQVHw5bpYDcycq6ZqqhPmwWyrngejQsFh
HN/XR4eRor5s+cGgfdd7CtshdI0ll8YtwUYR6UkhATcUkIT2/fBrJP83JN/Xb9TRJJ7P74cR9F7h
SJ4CGq5yqI7t8mZfLvSSqmsMalJX8EQlE1WbXNKH2NT1YigzcDLv99/k1Y7prgekwxgtaSSp09k8
qtXM5cHSub/wDX8A8VgMw7TrUnJ834uYvDwytp6KQBhzLWej9eWm+J9B1aQZh8Tljn1ODFxDl0Re
6AodMMN/GN/1HcP/2aCWrNYCPzcbvfDy+A3/KsZPEDZdS0y+XJnr350lTO3cqs51y8SF5Gac/PUV
N2Uqx5iMcPsZUPzBLyqGe4+7YLap1k+AvHJUaJ+w3RR7r0tfxcYYLFZEBK04ol3jutKDQmS2SZyo
YryU8FnXKgqPSbDEvmYd+aJi5qCmmj5hObqzlVO6JDvYmNqydkdREumayVr/fmTMEm3K8jOovVGK
FGMtmdVZnVyF5ydGwXvc+l4rAEKmlEDNuxS/67gxVBSk4CIRdAPCUetWfIu37g2dTmpmwFwdk5w5
h1vsc3Pe+Yr1FOGCzy94LWfFvsIlBGguv3zvusotGnEql27abMvPOncTn7FQlPMsPNGD8lqMG32n
l2TXKy91iBxd0e72rbaKz5Aoa1hQMWOZ89F8C6w/PNjs3krz7amh3Bksdpfpd8QellXzjYoPaNZu
jKvxt6vhk4MdhAm2gYcG/UHKoP8Jron7Kc4I+Fu6JG/+g/D7UMcWXvRXtsGLT14t2eDm+0FXuwdc
HsT94KdQQc9AkwaqmMwvncBdXI4L76QBDALCTQHaZ8YrflC2qX/6/rtsLl3rN1FZyPVBkREdiCjk
G9kED5/1XJFDSq+lIwpoO1ir35+Lwnvl+apZLUXlDMr8eBJRz4JBzNd0aMH1VVOup3tgSrFtomHu
lSTiDN71wnyXCmrrb+FcglWpQYi+N7BANb8kLR/q21T4WT+BOlXTQg4/ALQVabgstOgw3jvw89ie
qxLRcDWaYDovX1O7rt75SFc0WtSgC7rT+c+rfB5MMdCQVOX657RCTN+rNUo8waMB5cOYdBC5dYv/
N36zmL4ADuL07+I5AQs64gTyuiDxImrX0zX2dYUItW8dbMjR6CpiT9Bl2KmXtsWS/wvFH/8w8gXR
FTXbaA6/1o2X3DUQhsdzZM2F2KIYmv+o+zPjLw7HGjf8UiP60QT/CdiQn78qrmK8pYSPhG3N1lDX
TBk+Jq005Q1PVBZ1141CEvM5ISo20c49gVok5n1etyb4n1e3zFDILPNYX2YyP4hr2m89KjRCU7IR
RfWmm6asVKVslcXXpD1z+7uRJppJj90I7bUSqeTGN5l+xq9rTCOmY7IKyuYxTfh+KKdlEQ5/P2QK
DeKn4fpCRxlrVqI3bSlA2vzl6iYeoH8fXptxTTtTkDZGyAPbU4BAh5cGwE4pnGzWpnNykqYrXcDt
hidxQt+fvvHxTbsXtoB4pjwVXbeAsTyvDAohcpMwNlHP2mvsSzga/MxEVoGRAX5GSRnXbyqkqgwJ
z7jO6XdUMD2Bbr62vlGRye8rp8e52ytnCJEVKStxjOQ7f+Qud3T1jOBjNUSDsxkijEnjbGcoBUIP
bLveaSTGraBE5yqic/O4+dobW8KqzRXmYVOM/g9HiJ++2tn0kxr+8YPEvjOY6wGo3DTTu4XfvBF8
WJiKpaE11vnHi85uO2BTrhNblQwvw4LIGVgSMsDUDLJjkyVcYsycbY36AIqez/KMor0iwscE+xKS
o/O3GimPtrGaJYc8nfsgi/rzXGHbCulg8uAIFtC3h95zg5+ZwhgOcJeLBf+mMnaeGcfTRccFIZ7/
ia9HZQu6d3uB/nfZ+VuKZ5eiqjwVinGiguw0iHTIH5CkupHZ3fuvPW/SHSooqsXtWaObs6I3bdgF
SiY7r8TzfGpSHsT8mO7x5t3MPs42wOYrsT5BPMqu1eBKuxwMlQx7XTdSrW6qgOaeETSithGNUoQi
d0/hSF1VU19T+2VfTZd7afCPx8foG38LFq6+CV41CEWyQhPYoevBeVJDxliUunyvtdbgUG3TdFVL
3Uzc4CaHxzXdsYodq/7JdCNQg+dm0LcBRqXnLLMEbCCcef2hENBWBekNSow820rFg7DCrHxYdsjq
RhFnCZ2J+HliFEVZ7UXxrLtILzbPEK9SDBmWmzoaen4CO8Eb9bB9sYnGIojFr5QyAbBGmTESoTK+
iPGpTLF2+7XnC0Ge6BhkPuoPQnoTjGFWG/HlggboGQF5D4L44ApzotMeXPY4kUdnDHaKNX1QlG/m
E6HiLpLwWnmoFxfN07dREFVkMvj1eBSQMwF5OXK+Ol4Lpcz3ztadyl8XXKJPodyjYm9pwU88I7DG
hL6P3F94xF2luAdVc4YG4x0jsPnVDDDsKKrgF/WtiglCnzVnmSxtRgXp1d8nSdHN5Nzm0tS6D/7f
dNHftivCezbuGaFjgZzYoD88wNCxXU+twFc3D0UWimOY3BRsoeod16uB6HRQMfNMCJeWgCU/ZfgG
KWLh3BrZPAK/RcwyIyjZaxNUaoDrt5eNLx23/t84UhIqAB4+26WT5p6ETvu/rwpyFxk3FpakP2yr
EzAD8He0h9QWIyu9PJxsZi5Za9ZDeMJMFUb2+RhVgeB7T5i9wMISx3MBK04z3hLFuro8+WclPyf9
YiRRjUIYV9lbLS3jnjFfvpHeQDHeaBLvv/HyF+JHHb8eWF22CHf0ivJbuacXKusfJA4vponcTUkn
kqsCZ900rT1Iy/SCykQsgNGJFWB9RIYVZC/FM7KhG4yYe057ON7Pd5jv+YoZZwu99yOcKKnuM6WK
FZhHL1ShehXLH6DtWmmEt7XdK3+4JtzofvzrOoBlV73PuSq/uxJWc5cyIxF4xR65HOpVdmltYZ5R
C4EyW97e7d0WLEcDGemU/B0lPT2e+hRn798h3HYe3NUrW79yg6fDx/NMQja0++pWOtSPtKIbgjmR
eU7J2aL64d8giGJ5v1epWOiMoMGN2gpYd4dm/Pj5jCUDBEr76tuanDZrh9lctZLO2AlNk4zDmFDV
thhi8MPIxT+g0eqJK2DRVx7a04gEf8kF0lbpDnNEh1C8FCVI3h/w6NIwE7uXXzPtV5B5lAhGWMPT
DKELKgX3hr79030AA/tCqfJ3isT4KAqe0BlE1Wo3U7TynMC0YIwYO9ESdbT7Xo8PPoLXDPqwLxu/
Jdi3Fn9oc87cMjLrG90+Ie0yzrcPjSyaU2N46y0+ke+ynWoO3twVeE700jA9V41POJxE48JAE1SO
LRoslArP7Y5ZUC79xB0UbmlozlU+8pox4jwpajq3THV/56xqh7JCVD9GGwqSrRudHoCXw2I0AHmD
gyAtKFakoIs+2aIqO7cK0tve9ylM4WPrdyeoUQiPXkUubc3R/1KThj9/jRvvL/e6BS9XFNr8cX+s
k16kzVyuiI3fY+jsngni1DgYo09yZfmYiUD1AeWeXdpK/A+jH4g1JW0l+/1/vcGH/t332MIHtBOi
yL/KknxcQf7unyyH7LhuuuXMxVUZKAK3T+Hl7r3ydQJ7iioXnXuyWI+aBKbHarncAxWU7P1mtAVA
dDzyAt1SkR7rixEfTiUY0FTnF3Pvl3LtxwI4coGlSZK6+3GWqlm3lweQxg98ljPgRgHWxVpUCoOR
FmZlb5/DwMgZs10rXw8Bczf5UJ1F0d6awah7QYSIThHgobkGF83wJyGAHnQtl2eAN0FnvLmdoBg7
mlS1YmI33uKkcEMZAMieilJNih4v4/ttcEkQTy5/HX1H7JEfgG0Yof4WAok+/Zc2gUJiDb/N245k
ro5mwSedRkxULzq0fZuJQE8zbooovzo0UXGWU2HzByWYbNKFuzMI3KaXsp1r+CtcAzg29jgg5AcH
sA8YYMu4IhelLodpH10yEOLdDJc5O4iRuIBnQLLYdSqKU2ChHT7X1kpqXQLoUgPALwb6KaOP4pW/
iEwCGhleAnkbQs06Tfx42ywDvH95LoHnncW+7rLIK1394NX/IKwN60mDZ60fMG9eJcSGexL41BHX
MrCajXpovV4d2uxDdgiW/R1MNKeFwcnMk3YaakzxEXszZuxz40jJgSErdGEJUZbX44nEmnEL1qUC
Q/IuArpiVM1Fvvc02sVnQ84ZoMVJl24K7Z2rgCcGtu84byLUpoE6eNZodyZHSP2H/wy3RN+c1wEz
8jpyIar988JV75zdO9x/oklj01Zg2iD4OHCEX9iH4q74DvJg+fgj8a65/z5SgXgGUm1RgRInsDUX
yQtQzvQKqDIx9jgUTXB49ioz4pxSe1neciVREiWdmO7cemmfHVp14PeqU3mYVbnSMJYrraZH9E05
ctSo6kYQrVYQQMH3TsS/k4+Y+1U9XGoSmsmF1ONJd96Va7FxmbqpJnS1RrO/WSeiHhtnkzNcVJGE
EZGVzpS+Qb72llz41oK7nz37dFDCnYljC2AyhmtTaQzXlwgrdOMogiargad1Wl1zabN93d4ZPxDI
a7eyj7S8/0HqS0bsruuVrv6UmW3OphHhsYrpZXDZolBjyFqakJkD3Bu+SODqXeRAATbeit9PLqWR
a23NggR8L7k7BtQ63LuRx61+z8AYJznOtAAl11hGNo2W/NyerDLJmt08d5RY2dUciN8tSivrg6ft
DO7yRLSuJnSi4kiYfsjeMu5hSHmbAKUnW3FLz926NRjAqsrN5RmAM4fdIrbiytkjmL97L5eQXn1J
2MdWopE2IbC3Q7bzctG683cCEhKXOeUXPU9WqWGrW9xLVDOkIPL1r3PAIAYeDv9Ck5WRqgNSEyZu
l9PTkIdYQelo63NSCI9B/b/TEdsg64TmhwqU9dnnOdiTYtSDnXpeFkAjyRLJ8yNLPT3ZJwXcxZyD
Mpv/yEhNS6DQ4UhY7WFYD8kTBAQ7q0aMPNuP3PZxZ8QpCKxf0b1h+b3Pl6qqqdPHN1GpY3btAZs5
sjGgJI1mMbWxLIepET/AKPrSge3HGwBq1P0TArbqNcaPGBvtEWJbvm+rN2Be6P4HOyf+0qgtnRME
ounQRs96XD65TTNdkH/llJ7vIHf/sAfhS3X1LqZPJ6KegK416f7BXmTG/KjD53rncTVgk6pUPA/V
/bjR0hf3nSp9vvq/aJ5FgDLYHatbIIVkAx5lPHs6AhDMEc78+rgQBJ7wFB9M/RBHgZihIE9iKn9D
FrsKdklM+FA5aQUO3fSCN56hY4wE23DSUSWzAB151blczi0VMwfi6ntvmnnYyMv4dOI9HB3Om+Be
KfZVcWcM4tYtRwmBawgIJPzEYT3nEc8bSSqM8Fj4Zqi/3EWQ4X8LbHHG1ZEfiYIoPB5YceVYTCe5
9f2Pj5ZlfMfMtip3aVVv3Qos9Qniy3yeqK0x82NzhiFgT9ywYriVRVc+FC94LEWn7YP3FRUI9T70
Z6UpVdC+WpM3jYz0/HJCUT46xAo7ExVoWvalYE8PXSkSxsBCux7Fj/g/vQt9UT695RYlFqRuSRxJ
v2pxOJZvm4dGIQFs5B/63F+VT/2n0I7CPcanI1wSzFKqDN402YVsltZA26rLctT8v/QAonnJ6PeB
pLrIgYg4eVBBOiXgvJlqstoH3m+/LSe/EVogt2tE28RSdIY0918bDBtaYEw1dQ+j65btFm1TEFg6
wwzRHSLylteMovZRlm5rCnSMnF80Ik0B52Qku2eLUqmB8YsQkmYOHzKTHbh6mS4Sh1GrlCE5bXAm
jX8pQPs439fisJ/sEkQUzqM9H+fOH4IoT1ZHLNM+EsACoY9JYhrs0UqLtEG/mozHuRyu9E5k4XOq
hAN1E5qHXydY8w1bucSw4WzdTq2itRG+I9KeNNThb2LrcgdlzCBMJkcginIvPBAnwm2ohIHjO9pW
jgRXVD/WSuL/R4hqqyE/gFFXHNdZ0AtfvyvVOdLk2vxibBc56MmDlKra0P7VqRFgKUs7Mkqmqv5l
z8QK2Bjj7GGqGNr8hLkO7WBDgdqOs4Ip1oKYTHXh04tjQRX63ALtO5sTNlnY11Hc1OlDs56WvvFo
vle05OCV6qbhCIF2CIac4DK6hiMxdnQxMzFA/m4My2kheGXEEzESSHzHVVUBBgl5suraEagSqmxl
nBUvNXIz9sQE+NcOFsEFW/Ywm1r4lOW2s6tYhqOaqowAqAqndd0SuY3trdplm7Q+KCcEPz6DGcgO
LMylkdCopZ1lNAMsSe6c+HtkaM5O2lvs7SGGsmyKS9cyLeQbSj38q/lcYz05b7X81ps5xBxcBs1X
80MH+uERElDcpsR7QheS1SuVFiu5wIF/prmUF5cQ7mAf7hu90F4MmDxDj6bIQmyuz4wW9pq2nCyc
D+naHjPaYgIoxtwujI1T18C2dQXVzXKDDg3MTcD4xPJXkrq/eGYyTe1QY1Plv2+rRr5BRbDzu4Rn
+1/S/9jYzEuzbtj57DqzTA5oTTZXXxcuJJRtmql2Ff9+65xI2Nd0ef1olt5gWWx8EuQIFPqixc4t
nkdT8IDh7j/q1u33eWQofaL06vZCCh7Jjybuc+CdeS2JhXpjFUoByR/RLfHUjWYYEoobStTzcUvC
AOUOvEUj4qb7iIqQ0eCNziisHw6jN9zSVbhJTWs5BIyHvvqkU8FdY5uT9yDSFdWfBmqkAU1y52qH
QBUESIVaP7WIea0GzbxbeTKnOWWRAjrNis9Mq8Ol38hdWaRGA/eiZL/7eoHETD/JOIfQUgudpYJL
Zpn1uqf8G0nR03UZsQ13xOJFXWr6ZLtuNiLvE/wLNRcHysckPtNz0cLMo+7ZB1h6oyM2PuMbS9QY
Wgl41J/6T9KF5x0woxlQmV2XBVUePWWJmQ2SBO/LP3YUt5XQ/T7oewbRsxy/FCAcae21uh0FtMMb
RcZv5XGsZyffhlu8emKwky45iIK47YS8+ZqDoquG0DNHmyUAHL/fd9tzDUUdSgq90V5MlkOyi8LO
6SI68X3JD4kqCJRCzp6h0SdyBte9hjaOGi8ejU+7ct8qLt8lMSnJIhAtmz0Wn5UOpF9InWWlVZeN
Ru3IRHpb1untwnayJgpYXIZiqwZAmh4bMpw5Ssxp4wUgscbqjLsyGbwoHi4p9lTPJn/wiPFsxvCg
XPVYe8U2mkzC0Rlc7b8unkPb282t10YBwQU8P6lXY7Q3fGYA9foHry2VWd2c1OyEtknS1Kk6Fmtj
zKDViENjHo9a2Md39zfuunV5Ypa5G3MlH+z0QCcqJ7K34IP/6vnqSb7AqT8ZP2cY2csH+vK9x+BO
xdMCnIvgJxqecLY5fyIM9fST0d74Ow1bKSoPuth6nHmjGcXdD3cjHnpoR49Fa6BQlVa8rbg3HjYm
ZVGy4M/KCn7UelYxs2OydgDIDOWIMM3KEMzgB1uG0EyUEjUBTJWrpBiz3EfxBp25A5+JJ5khjsBq
6b0XsaW1Qtfo3Im4YkFcDcRMheQc0X/ftX6vuvqRmczH2GYJWxcoJ0EaOlJa3KtO5S1zA1gRYY7w
zNBw/3nA2qMIDPHcH8Ol+qM3K4JE7++7r5NhS297XJXb0w+zFTOlE9jhEx7Y89mT9qjjR9y6wGZ3
cWYTWINft+6o+UTlFFtHKN/AISUY1V4b5F556XvXn5L40VpNRagrmB170555GvaSgNnDMOsbMQrh
uRDr14ql0gCYHcZN7RDwBdw7AH3X0laDua5NWUIVtklffhFyKSdX9M2RSQAKPTEJWIGIjVvhO9QY
V6z1wQOPoGAspz3btyT8Ga4+o2/uTb8EX5hgvfF2xGbMUOwc7stVyEn+eS5Sv73/HTz/uLucF8xf
8/9U2kWzTSqk0t4bySzPGyPkHRfYcj/HTDiOdhfTh8ZyCcJXA32dY1T1gxM6vXPBIrHBa1Uorqmt
Kdl8JycK/FTKuRudpYmOxsW/jLCIQeUSAQlJ3WKHW6oyXolNLvMNBrX2+lheMJ5HiBXw9JZFKzy4
TD8khDUHAfz7OeMBExYyNlo9kMiAWso3Y4qIxuTtA7At75lTMZ2XO2uwXym5gUrSnsxcM6V4iYBE
Kp7L4pn+S+rPklFx7JSPSndlHkGk82kxmIXBUnV62Y61veEjOPBy4zMcX2JrrksRsPNFJH4v6gdA
VsVsl1zRZjdlEzLoOv13PlEfJx1kIgga8i/fpzRsMgzV4556jMNDWuBYzkVUWQ/aKaDRcl1ELvvX
/8uH5SMhFMi6SV9rRrTl44uukzvXlnyYkSOFHPnK+VbdvPN9VDtxNs+VzklufiedDejplvpDOr07
l5CKVs+fHBzhmWgZx9rzmnQ4zzuyXFuRkNeraHrk5Pr64Ni0gJ5ibVV4RwQHEUEjke+93S2zo2j8
y2oY+7/I1qX9mhsn7zC0x6EalOqFIgHTyVEFA5ivirWdQAw2Bhp4D4VpC8sCz2ltc3Dn8Kdqnk2t
QBdEkKCFGpG5xLP/cpDQpVSnlvLTQTp25490A15G5DZKYNjA5Ql4Jey3YYsbtackZDnqDqYJjK6A
FE9QgF9paIciB3046WtYMc77EOpOY1MFzSntSJTGE0eiWbq2iNCAI1Lz6BNXi4i39+SFKmJmBlXv
TTVdgfYkOB5ZjLLaX/WQXYNvjsQ41bfHMwExz7GNLfNbEUg4dpb/uA2xs69XEv8ctANFusxcYO+O
tYp8lhpLPiNkignx7W6MXFonRdc3kOgwOMhjU5hH/MhhNibnAsn7gUMn8Uze/jF6srIqiiR02m0v
rjebO+dZgafnLmmMpbrTgOlzawCY0H9mGLBgjEhk42W4x2YqzIVDCZ2a224v9hbtog/ebhQB0GZs
YKdjBJCPIKYAcYgk7gIXb33IBJhKhvEBUeZsfW6/i9/uNkiNrvvxNKbRTpnOwjnp/no4T3/etzOd
Bd5kyUWbgtij40XCw9XbEH3QcG/j/3B+2cbf9iPVRxkDSKo+qFlQZoZBvpi8OsmPwRA0pZR5xog6
DVa9rvNtuI4a3ffAhM6bzpmiHfjQ9MjbE3MehOSrZysUYhpuUF90l/iES7NFTHjbPsMz9VruyH9D
+jsAkD+zwua48r1LQkEf5GaoMY2/5dZYfB/Y1asG/yAkbhFhMlsBhYcfnnc91LMSufuAuzVH1JIA
m+4SI+05htAXiZSfVG5IUajy4hMYvdSZOaichhis9o9YqBdhAlvldxeJKCA7aJbj2PItwba4VNru
yebX+bPsJwQhalhYPruWuU7A1yR8MQ8nP+2thADeDINl5CjDBL94Kb1SooOqp2eFzeOobuI9xn6e
yc4WDPeAZjtUnaja8EimesCEYcwiNLj3p8fwXVi0RFkMyBeVHSamvUt78CLW/Ar77Cglim3cvnw8
eymHKSd3jaYYAj6Jj1L5TOmB+1GGwZBtp3/4mIrpkYfcasdHV8F7S63Wn0r3bzBHisrqdP4bz/K4
MjA7hk5nv9NJcgqHtrNFrT/cP4DZu8d2o8tM/rlfZl3t3t0PHK71jwL6neQ7cgDTXm8ILac+1m6A
9Ovhn1e29RY4OOCw/jVXsO4xrK37X5MsPZcs5ZxR09PGZHow76n0ddJUIPXpE/BAvefR/PsESeV8
XnK7E4sN0jRwJLIOhAHNWY3qAPVFNWX3xhqi4wtlwHwVmdAbQNrLB1O0ciAr/YJDJuqoXhuVK+cB
Mm05TbgISWD0hQaMMLatqH8RJKveOiqlWt4HaGFg9fjJmoAHJUvCjPdIsqgswjJIX2CDL12DJR8/
3v9EB4bD3gQh81oxQGxVGMuOFtg3AGbRA7XT1o/q4nOsuIf2n+4vL5DZLYHDeyVug5GMbkHvLU4j
u8x8RfLMQGtPqptlL/Lck+4QZj/F6BDBVsrH+XwjTQ6XHv+xVumoKT0w1TfYhDec7AvAIOSkGqmE
+eapkUuTdBIeiRolxWgCDHZHLfcU240TyUl1ByuQqMMIY6HR9pdtNL0vpaSVkZwUn2fRmKZdkR+3
QMa00DcmNium5nP9bQq6WuuO6/PQcy9BZVPwEekOFMh6pxJWBTVhPzB/Vw2p3ajQoq/98wuXT1C0
Uth34KljBZdWLi9i68AnqXlcurP3D2C2CvAchNNKPwii5TV/dTEI3DJ6bU/JEzd39R7tsUmZjLPw
08MGLeRuNAqR46D/c3FXoAPtro6EAlP/Kq1xozNMDFtsQKyV05yVFI0DTlVR4Wldy3UGkJDBFtU5
GMCwFiu7xtXJ97tUno5skGk9M8fcJWYcJwQgvHipOEobeG6v/864e+eJ25WMhSpnpodGlTs1h5U2
kOna0INX3O8XkJYmVonCv8L4jnD0dd1h03b7XAaMGhlCkdjO1K2IFdni8c7k3rZAxz9r6bCwK8X1
PNKoZwD8d/zsTSvvclGVd14bRBJ7PVseyPNymM8CA49NbE8ReEXDjcqMDCaUkyj31DF1/JKY8SbK
S5je7FD+jCiEZMEOirllRROfjMZieXWAhyZHa/1ydcblKOLdpscoUrHkq0bnFCTaJOKabyTGr7E2
HlOqT/7cYeuLtui64X6mR7ST5MrBwRWTETWYooMzEg8FWcVUGYYWvh8Hlb3rl7xhZWF9tR21ZG2F
oRZj6XcxBc7cL/Svg0ml6URDbzIpENBcVl7H+/iCk1Kys7MEi6zR5x2/dUG+Wz9qcFeqzmsuDi8A
w2cwddyzeoCdDq2owpZpTGOw5JnSCeWmzHzrTiWpE73yn8LnhRTB4DM3L1ZG3OO8AtdbeBvZebD/
g1ac2vcm/F5WG3tMOOdHKHXd5a9e/v4M0/UesTUJ36iO0e9pMx2rCJe9QtX0sKsDiZPzgAfFxSlr
qbGC6iNrGzcgBt+VDAz4diR4kJkCpnakfKif4AXJhWGWkYdp4I6OHFif7h7bSQZAk+6M/wCi1hZA
wtekP4gJifJ3Ci20rqf/K1h1YRF3HJ+F6HSQ6VgOF9DUF7c7utzu/NZkC8Sja7UPXD8S6g2pTAjA
jsY8p5+McaOEKvGJ4evoAYFfQP1MQzxZr621gLbFbOhM7V+GBTh6o8Xxi9ER0Rn59aFZJIz4JYcn
NXQyo3f5qXOrGEEQsfp/qplp6AZSO3WCwnQztV+e89EAkPZj3qwlI7EDSXF+Wxxo5saLHYza9mwn
R975QN8bmiP0ApYs2LErIspFdigT9v0HkvCOTYYrB6F2AqMepDgvQr6JmjYeIOZgGGdsNvWPFVuE
Hj2BmtNsfRPexyd7720wMP76po0f2Z2hmFDjTfMYCszkekCSJyQYbiFbjBkeaaVgJd0/NMnN8e6f
8+s/Is7aBXryYW2tQ3kFrq5505gcLr3CKEK02RsmWP44WlhtGkFH+mhJFt4vOgT5wDEgJw96SdEz
PNJ7jDtzCNfjPI3J8q2C/ZqA3H75rJ4m3igR6cOxyqG8bELvOJDNIKCHbRxg5gNG+MaN5HtB17ti
Om1Xj2z2Ju+8v1X5FFQWt0D0R3HT2t7YxkoCoIFs7ErN6JuVoXP+zc6mED8ZHh4RecRMVJM3f3le
/UtqU7MfjdVbT1uDKCKjrTIcN9uXN3THZL/tSIJd+OpNMaDSlEZOWS2CJa22rCGp3FyrtOeph+Go
9FAM9HxgekCGfLZxdyHEoiF0aKAoMaVmVilj8tdwPtnX6Q+C1lAqBGO3S8f3ihzJDkdMg7IIjKSi
rzDuUFTu1rASdmmtfqZJ8KZPTPWOAxQu1Inrry7M7TaNXONVj1RlE3UVvIoXlw5ZwFbzP4Zk2TBX
+ZZdEDZm8aF9ZfHRX+G3QC9GUo3SA9d6ZHlQYA17RWFNlXZQaPzKzWMa0kRgEngbI2VPBc1v7Z4U
YGQZ99ZFQSs8K5bH666t2fdHQDS1p63U6sFwev+InUyiUDHpzeJKrmKAfOJubXowHJxISA82aC0J
DkDsduIJ/NZVOZpeoCsMBbfFvda5oAJf0ItvH6A0qmdXMZheGT4kygt2rjqUxVlzCDvVytWEDUiW
+LBLRfYm5OqMUsgxKfbi+sHANlMqDSNwsSrSPyc9lqa7S4mdcrilYLt/UYD1fFWaL35MCM+YXAGP
RE5qi5nMw7aYOZc20sL5YKd08Xzvwh+2OelHkjc24mJFapAdimagRJxi63nsOAOLeQWUaZTIA5rM
RxMHZcJUdrc5+0v6xuYUm7oQN//BnM6dQT3FlYRwyK28bm+JmNmVQyl3d8vGLv2pL8Z2jYm5knOt
gLdFzOedVNPnp+LV5xkYCH6AxciK3I0CipkxOYR+ixGFZTjUl/3APKFB6My2c5cpTp9Wup1WVEtK
bRt7GRZ5DmY6pdYzKZ6sWKvzf24BT9n0l4dEsoPLjfzzip7rMqTkD7LP8+I6QdKgS2A38eJlJhDE
e+oKwcJHKac4NTVa3J6CfwAMD3grTpZNKwLSwdRXoQrYdqlGiihO/j3OPZZYOD6S0KuKdJlrR0Mk
JizplzZMXYmmyJ6VlMEH9hRmgIwC8Y8xBuCQDEVc7SccsWa3jSk9MOyT+BsZHGWB2juER7iihApn
5K/QpYAQZo8hMufNQMzl8ZqAJ9OaHFT7yYf0Osmzu3vMSPbnQeMbxn2JKaTwIiw5ZmciPXCAUvMb
RN2EgcpSzomcdla7jkXn34e8siaM4X1NN0qGaDQxBNSkrnw2yD+tMpt1yiBjBUJXgFEGbTHaNYXS
5koMHNx0vrhTmHxauhU+AwM5PV5dqslqlW9NoLH1pnVjo09+8wtDfBflqZNylXAdTp1oQog2wtjW
2HklCb6IUeE2ToihfgjFmuJVd8CI2QJrfDQLONel5J8kok8fOzsg9tRYXjYOMKYOnrVkLSnmlBwP
vsqUBCGLCBS31sv3yhpQwgpaOWf93ZbEnvtoiTl1r84eYxhwD+qbBhu6lkn+GASdRLFLDknoOdqy
F15gSWMicEi1xk2L2pOfH4uMUXPpp5QZqJZTCu/Xyk18wICDrt+Bgg4FvJeCeRh+jhFFSNh+/zR1
NEI+SPY/pHI4SFwIuUmLQaC8mHgGaepIr1mx4I+a+jEfleGmR3YlpZXo1l7EsLmnwMqRJeg5Qt0o
wIvTazFWRV2cxe6goUqbVW/VLNbkNLVLmhJBzEKjofVafOpP/1y041BToGzgoM0HR+2qwdQtHIle
8jospACpSDT5uQlZpqRQpAuZcOzULhkwVRyJojlZnPb0nevm5BZdSQoasFLXo+NSxsQzmjcPUt3v
zXYHpwSKJJQyvRWLoueXp1n+EjCIZIGE9gZUcidB8mGmmR479h7tlGpFzPeEXFPjyK/3LDT9SHx1
CwS2y5qg6nIidvTvlkl8rNvY4mFBW+oFd126X3DdyjzNMF2XD8+Yj84OC9TsVyZZnZ1qlj+If4Mp
EvEeHZkc4dCtRhbt/HRjp4DbEgU3C5fKwtPBRII3jZpWNSFMkRooa7E7yR7cquP/N1F48eaiWNhK
y+rEhJBv3aziga7sqvoKgCokvuuG2EMMQj8XsCwpwORI7enqSL44/3oi40Ctfd5hreuy9AUEpb2g
yecYIqyLWmshAh9WTfVwWeKzDeyTvlhIP9WO5I9BOIBJ2UaL5zBnIp2k9Uks4pdTyGSDY12Vdqvc
e8WpkL+36jIwW+gK94QK81MVT4tqjUNdvj+96KY83yy7RpMSE9Vx/XAua1+Xmq84LPfG7kIt91T/
8u9CRs+I85hz5qdY4Yy+EoX8NrZbV0A1Y4CxcqM7qqFlgntbCrz4IKvUmtyyc24TOQtTu/XZK0gG
DWq6G4R3NLNUxIPx7RA3Ebp+b1ar3smFmSoITV4T1pzECbkY6LqofoacpGl9bq0KQbk/PqCoq1DI
pxivaSa/WICItbrVOPmY+f6eajLnK8CrwTnz1086vvxc48mbNNGFBUeTsp+C56JhIKosFpMjWD97
Omh3mnmDUkF9F5EDzquMHP5W3kBkEQuWx4kNn2rHTNZUf2j59VuHI7hb3LhdA9zExI1yoMbuUliX
/CXOe+J79D7FM9640JhNplqGi4oBtFqhMSyBXkRFwPn7toRFmTUjE8yM9z99QvXdeBGiBTTd+boI
KvOPK160wcMfm/4gi3Q2jrW9IlyAphYUOSwUYg0iDdHPXNwcvcFwSvMFDgZnaPzVXt8DdJFaQBeo
nl3bTttoaoTVHnmbDYmZlLoB6D3MGxiXpyRgSoCDRoUnF5XA3o2d8R+Hj9/Ah7WrV7HHOaD3XRXC
94Q7REQ0KlDkUNRM8dVkGNDtHwDOU8KmKt9t2tEhUnRe4LVbRussN6kWxsVPXwrkjE3YG8/WsLhu
caUIGpMlVYP7I/lBrtsR9ZEIUwaiKhSYDkW/BR48TFeIaZV/rqB6hmI4QH1N9gz4QsPi9F8qORt8
4n1MyFMWpCNNrdbH09vXrAtIDk011lYJQ+b/0ZD8HFQRrrq8Bt5r3QEw5SLEbu1owK5HunyYPtxa
rKDsV0vLZDNZPsd3HXMm/eArkrXZHaoaiXd5DCOQJ+dRVj0fl+qXNq/Nwqt9v/NTfJlsiN91gUa8
EQEGZlycDjQyd+DNK/JYdRypWoSaBsYAyp2qU3dQDGH4EbsfD9wFBBdWSrG4oS/lmTmXtdNpiXDk
M5VL16mqX8FcdxF81IgEjNJ6h1U4UZh6uYxkIuAimeEwd7UUqlOSjYjehnsjoBHMn7R67PBBB99C
R6mEgCyJYs8MWvjTFqyYZ/5xNZEHwt6umxnXGyuiJ7jLc2bY3HKRuLjCA4vut0MWAhaQM0IUDj5k
vz20BB45z+0jH9fUGgfcaZz37eCcdGrzaOiWE74GbjHfglRXcSIdvVT4Wh8cquEd88Wtp+Jinpr5
ALnuU0QPX9mAlMkA+5h1lCrGls0xPCvattP09T5Gf7Klz01CAZctd/oyoIhngzyw22jPaHmLFnsY
KLZ9i+fdvdY4b/bZwI5/eMArzr1hrufyfqXfthNvusi5MGkoGWWwD06WgFYkPheUvFWp9ghYtBOI
8O/xNkjO7KoyOtdKMo4qbVn953oAfbHP7TVHZtWqiuAE7hkBDBFDxSxsUnDhIyPAs57guTHc1ZXq
tWrYZw7a/C/AUAaRivm5eekmc+ftY0oJM6DkjQjCS2g7/P8mH+vbgJ5GI0xB3gpUOwN8cx0QqIjY
uewhWZdmYmAL/g7v+b5D9tVGWrvRjJO+QjtBc6kNiUoygOoNd6mWbeju7yCvhnCHVJK5U0bbQ+wl
JX8cygRPVVEibiZJ6GJnwGdIlHWiFbEXb8vSaFv5XbmAD9wUiRHt6CsHgeMuW0R02EX/7EgiIKQ2
/w2LqhuSJnmewaxQ/0+pkgEcTmn0JtXzhZdcjwkha9M5XZRR+m6LDHz4Q8/Fcu5AnF1CKUBJFvvU
oK7pUbzkjdlafK7MGMkCmeFL/YFv9UY4w/p4COeT/4A7bvC0BufYgfxEiLeTKNGQgOrzR9enMr+a
mJ9tvoquDmjNAjrPzRHM3ni6OZAPs2b7YMEgKgSdcJAtkzA7uf5CLPAwSNZtEYOuwyit1LRm7ukl
HJNddhC6gPkGtx0VSL09oQzToPiP6IAYy2Pje5n5s6gsjNexUV/hup8dx/xVk70ZkJaC1BAx7Sk2
i/cr+w0k8AhKQ6rq2nEXZf8Gco+1uXpp5UPGjnjjrkwriDImRjWf4NN27ka2cjZEH5UwDpuYVgx4
u4TL5wmnvEOBIKQna6CWjhS6NLNLODBE6K3oumHus/B6LcahWgiS9bmSGJ1zXyW80CHAVPFrHS6t
aLgQMgsNAkydHBrdap92GShaJy5OczwDS3TIgmyVMl0omCAqJqIlPKVFodYcOBsOpzROfB6gcHXt
xK/f1202PoTCBvuwttQNdGpd5Cn9HV8JjN3UJDu5pd93TG4qHOAQ8+w6XJqJmunerMIDYObcK0Wt
k62kXEMGfhDQ+z495wAyrhkM+AeEzrhRj3tM0Edj+BwQbCiY0pSUCRFA/jFd/LjWibX+UOWYitgN
H3XcsQ4YDeFYdcX1xx2xnKaB0DRi/ICXEjBYf5OhRzhD8bQbV1Xri2sE4hB/1Un/Qr6T27mmJt5y
EBUtJjWKcXONYa5leKwGfwDGcqGlzODbAhfc2zTPK+NlxvIOpdUPUJVKjelYVoOOesDZ810JnDQ/
i0xr02GYbjMB3fCCQkVh3QSdResVjbmy4/AnK0q9sChscmP5qZ3Q7Z3MKtOL684TZ5rHym/ly+97
8Mz4aqtF/rp68sAitRKaJvppAWZjn6xKRmpLet2KcY+WApW95PmeHWH59I/HDAJVelXRZjh4+nAU
CHKa2ft0jwLRNBMHKFF+Rc2OSq3NHLoBNlQJ/4iWVUw62kKeCGKQSgfe5accD84UXl29PiFSi4TJ
apGR5uxl/xaySGjpY0Q8Oj69JA0Djp7NxAu7KbJ+UElD/3sy+PrUf2bFgySimti7YTv6KHdfO4nl
AV8Zdomh5HlhFaGln8Q9IaLdn4cRPz3uTMt6q48B1R3i11IyeAn842fnTPtDnMRVZJfZXUuBpNzZ
CuIgJ9oSxe84vEokyKyr3AwiWF18wGdsYuX9LHZaY9dmwWgze6INk+2eH3adfVEjJ1SL+QJWkPf0
vk26H1HFvZKu7bb3YcEw/9S5tAKg7pu/nzJkHFx53+cWeGMS4238m0+g0lVhrqUNA4kVdtcRBP0W
uVbdS8QTi9C2unB1o+cghEQC7sEZllPT0MYzBASGQXXR1EJkSEJlqeqvwpT6ozgaoxfD1YtSAOge
MYFkDm6ZEail12zD+i1H5j7nmxEJ8isco+ZNoDTCETUuAUkCZUN1g9gSeDRvGe8Lfq1KnV+pJXPU
tw8v35kKhXDbF03iHL0sx9wbTgnHBCt6AzUtrfW1583w/m538mTgrsHbxNJuTYy7+S/5w/unZmKV
8G7ucjkoGB+puj7VJdGYOFz6n+ksIiDRZdof+IFr0QF/O+IptDfNvVg7GkPiZUt7cOAC4kTqiuhs
2A+S777OLvWNSY2eU+qxl2akP/xIqN3Wy0VITSu/I55uibEMBXzzysxqQti/Kt+FsaohUSj5YDBT
fd/d0xt15tdLzBp4qWwFuB9qf6nYgFFJI6q3jGFe+KdwrRCJ+Z9QQWGhan/YQUQ711IZsbZmNELE
Vn6DweyBER9UL++4kKP/X51v2V9lWCr1neUeVkRqfeqB0H241RBSUMxRV+HWph7+oX24aSSCo/Jz
iNjsy4kfB6MsNxIUvqyssJIKrIw5z7l189H4WPWlTabbMljJS/L/xaHebXZ1PL7xCajxIS4FpOkt
cRxZgYwYjqrTN6e5gQdwD7MsUu6fzc2X/HKkOzMF3CZhot0WXPBY4ZpSY2nc7FAuvzBRQf25ml4q
u0ik7cWx1O58eLHIy2BrySoKLRuB2aGYIOtKXaM8T37RMVmf/P7aLs1IBhIz9JzSr6WQvrGixLVV
rQlU34sHglEZHIcDswkzqzhee8565INqAGWXqCuYz+iAJPwt1LI8EZhw/G+K5cVH1zUt7TXx1CdZ
FHHTWQv46ZSPZaBuP//n21NEV+QuCvLVM0Yz9Ki1lXs9KfodZBCuKz4jqMbOiSjmCZUILBvypylF
mVQNcyALfT12Di6t8A5FZeS6UGokS9l+/1Ewj655DnCUDujme0ibJ304CLs+zAe9Z9iKJ+7tSmOQ
T25id5T5dQzYbUQXZ7ToWOGhelpIJb+0NnticzRN2gJjq3mFvD+NS071LBshMPmIXvUAUSg8QWvI
idTeMJvSJDZ0r9hgcz8VbqYNqkpqz1JaLqb5Jdphs28ueyB3a7QVDMkpMuDTfezIgvb+CtAUTse/
EP2so78xW/HN62fFdYx0xadDTSPPdviRDRJ0B4/CIeIHbB3/1O0gHYdPFzEvK72Gn/6RmIIJst+v
k9xjnPaUOTCSC/tslMDc67PYan8Gwt7aYW4MF9UUVres5Ky11zC2AhuXzWIx0RnvVS/qVi6cExzp
yaLNZb6YMARReIpBDoCkjIp+Js3pfpZQX+TKCgNHnVL1ENLshtFKdn6LZ6IM0HlqyXooPiIiJeur
uOzhEpDd87z7MZZu0halnnraAWkgqgyb46yreAb51+KG7K4Vg7XaEiRT8/w7bPb+XhhKJAzCtdew
SfRepLxz543dCCe/6XH0z0XeTqUDaQJTs1wffUnIbSuf3BR9bnQdPyebiCMyupp6HMvAK/ZZ1j1n
PvZV4tY9nAhShYSDZTvBwZt9VscJCI/5ciKRrENLmuiHx9EKRfHw+aebJ5KMWVY+QhRtI5Y5IafU
VFlnxd8tpXjsYe12UX/Iluq1vjdvV2FCOR57vzPh5zX2k6fBYpMkWcl+6HZX9BQsjfX42sygB7Mf
EInk6w6Hdwe5OeEcZ8Ix4g+0plEDFdmmR5CF3GV4HJaWwU8cMX6LY6wCyOjBJRchymbScZxmkpkX
XmE2GWK7ah5p4IWeeF28KHwc9pvEWOLyAo0njGaZCM7xHh0Aj5aFLHHSUYe8ksZLRPKzw/SIUeCz
LgbRT+hWIxZ1eBFdmtaFuuaYTs1pomQxzlT1t6s3HQJY7Zl7eRTxvXUjRe6FKnn/RxMACoM+VAMR
iJEcyA+ZpcTWd4lVS6L08xWSQ7Mt26P3AFcG6GUdPtTpmpNCb1ZRqx+FWblb2A1bgVc068MSaOx7
H5NXurpJ92X/tTdsFOtqkt/G99Aya3v0uejOvsFX7T06b7CtJfWe/GBSmC6XInvixYMiesxK5Xem
w2BEa0ukGLm7kij9sAjcSjaGrfxSLhojVe/tjMPDCsrb07XWG1ABKuEf8FKtyl8qT8f69wGROFTD
GA66p3KNMbc9DLbyg5ns+Rx8TR/cyOLWlgAPegIHac9nss1rKq8wvst7/o52PTML4k3cZDsFImWU
Bq4WzlbykeUHTHsVrLq+8+LwcoTqwlamuzzmkoZyU/Fd6QBpbtxHrws6WSxRsR3hy1bFgxpAYYlh
S3GzkmilTzh0tr+o+Dj37L3mdlziM+Gf0JGPdBq3b8P1wPs7lhzCK02SY586rEA35yEEqpTN4Bji
VV4QvWdIcpQbL8orDGu4z9Q+v1YGCke9azVuGTndZRB0qt5qi+WQMwGNplfV8q+5Lkzn2cSAwvf0
B+QZ9Cffvwn8zLL2idYJ9TJQResH/rG5P0zDgqx1LntdTTpXulERHp+iz+FBvguKX9kuobLG/MIt
eO7JwG19vECPoHmdMZi3lKXgGRPxg9GbnLMLc8rYVUPqKY5LKEtDRvTZvFg6OutvKY2kHDPEvDSg
boogiLdmdkgMWxul9t387i9J1W44HoXKD0gYlX0Wo1lMCmRcc59FJcbYzovuUg5H8EDE92JYvmS3
5jWSgJdECk4lqclQecJ+1RmFnAPmmpaxxeEPLIdV++CZZabZEkkFyJN8fcgWubkUKq+PSVvQIZ9Y
Ly6OFhifHVtxIola9MHp/o106SLQyKu7uper7Plq2XiOOnaNnon2iiEd8Sxmf7VWMVt20V1QU6Hj
t4Fjz0kgsk+rKOqBkCHsO/ltwdo5+e5ryzwvcAufytTReLq8zoFCWeXNWbElN3o1jBmHZHJg6Zol
tcol03DUo1iNWSqzhOK+p0voa2CiJID5vPZnGEojWszsyBvV9Nn3SoIxrmfpSY7gQ+3+atYEzTYQ
MFRE+hz1oQN8O5szrt4WJT59LHdAbz9UOloOx40bUuryaLu4wJMmxl2ISi4izlnTBZkgeWIQoylz
QnMz2pFeGGeSAe4rCqjcyovHRRy0nZKvu6kYfCbn3da51xTusjeazccoN4A4piZ2hz/7qiujWtNu
WKUsLkaRkh73WyvIvVoVdGV/IIglzZulvhLlBFfsqaUdWa56nR1nlmdYv5YNUwePyp5200HllrmB
Io7uBS1YSq5rdDTWcE4knYWVMuql6HN4OwGaw4owBnzORfU2SAQNtAZcMG5/HyTDhTwI9sLlXWS9
sFJh8bFBet+0WgZgyilKgYT5FTt6ocgo7v/B0eXFM6BZntWvxzhfv9FKLPbIJd9svC3PN7UPjz0h
RShJJ6hAY2pkS3wYu4HRnGxKF4wjAhi52Oz6pRP/VuzMhkRAA58MluqxAdyUqg3ClP39KgRRjicc
u15rQs2ahOhZXStknOAG5ychbX0qRMC1HRMeRO4yv4XFUFsKyQBE5SqMhZg2wFGqO3qAa6kjV3IG
zOoVxusF1rdxmq7GY2CpgOdL/P0dmWPPwJ+i/eNyBvUeXPo+HI4ETAnN82Gyl617SqPei8D2yZLr
PtgXLEkAyBiRp1OTmSEn+YBSdNA2grMSZniBq6O1fc+JY2MBJGLhPhdPbibkTnGi8BkTAOII8HbG
F2MC+wUKWa4UdVdOd3z7ULc0yX7IF+hrch4zZ2J5pU3QsstVTT5IjR2npL/OIhTu6ZaawuN+I8Lt
nDhOinwZnaM4rxO6WFulwNQBVMnMf7ArECmjEOtrWvFNOnbwUsMMkJMuGQ8ELoPafS4lqXofLA6t
EJsrngzS0dXIRJXyx1NxvVXEUixWLSi0CpwILY/rrgPOzZIYZX7zIYJWwAX8v5PmSq3JH3YpwYsG
BjBA9C0+jArizlF+cdVLordUvsmLLjwMdWQibN/yq8kTcQ8a7hUa/pRZMybf+wc48oDmq7hENSht
MQaKKuBaWLskpIFk1L7ziMRKji1iQGa2l1Z813ssPPvXtsHpx0Z0RYCrN1dCBnosEdMbrUgoVH3n
XH0cMohbW/t7B/7CldeKFYlqdPOJxz1BUbzxdzgWZXbYz9vPL4GEoGXkZHcJ4/j3XBM5Y9EqmaPr
Rv71TcUBGiQjrRmUiDXiJenwxiYToUGZjYOZuiYnEkv1sBv4g+vlvDGigs6OSdq9su2TbDZpdUhB
eD+nliYQZR53pmYkBCVxQZVcQ+4uvyn15eVMpbQlD+SHg4ER14lHsP6wB6Tt8qPn41rJcP09T0cA
txEhW0K19xQoapICH5GtaIA8QSir5y4hmNhXhx8wTAgCoP4DN378SnPBC0weQmMv8r9WZnSwCPAf
u1W6blAzlxOGDpJWhMj/iW8T8VSojqiQyzEFyYK7eApDPbcxqFEIt4B5SZzBvDdnBWmU/3aZr3dF
OqaHypnVZVFTgj9/gvAj6o3sYOFEaoS96ue/mMo+PqW/INKAdaYIGZXZr2jZ5AEITm3TclDpGb4M
v1gyA+Bgu0LN2T0dj+9Bt2klhhef5tHvI27egulL++aiaSlSe+spURVAKmGNXZk5VkLQWgs+Vt1A
Iv3vK7mOQoczBJrjNKeMXFhP4SMWU9HnpbTEHeuSDEeZ41J0zD26P//l1IL+CJ36W2V8nZwbQi5A
cqEzvpFsiGIPln45fYbSxHEidgNpgJH12zCZE7GBjG2bNlZ+96RJxeItfM1Zk5QLRPqKFnYi72tw
Sg1QzJ7kcdTWxwHePyI4mSDkOIoWaJo2vQuROeaJzG2nZN32CjkHl2cXSds2rWMnZy1Cpc/mR3s7
vXJAiMQIR43MD4oI2613e3ewZhGdPPUobrPqkn8IGamLEKW9H43DeabJCkMEglrWTfrDYRWOCaEO
PxJ0+Bo73FgOmsh5CSMEDKdJQdt4KT7b0uBU9hSZ6Dr6FH0JhQaXrvt9vCjLKOcGnG2AwtP6XZSl
GoaEhk6KGMKb+OOiKxnwk3KZYDAliLwQ0m5dOC1fDP5i42O8n5icnNxE6CXZothxY2eqe4CD3fw9
kubtmTQVwL85xUQD0dJlZ6XYmVJox/G5VrqPTd9O02PI7tutRbGSiT7P7slPE+vx9ZWqcBZU5JKB
thbkJ/lRqqzRVlrDrU+CrywxgfoIsC6s825H3RyV1TbzfWwJhs88Dy6Yd9ftA+hU+j9QJLlAuY2f
A2XK3PTCoxUP1FsJuKuVIAeU9IByGJHIcfLVjtENh1Q0/4xOrQqmaYvSRJB+8Sy8g/WX2WnS1V3v
i1Nb1pAH0GdscqxeDyJhKxFes6Hlx9n3wlQAw448r6URUOX71AHCiMzNGNjs+nu1hIJ70Jnobo8P
tC+7yiTJTHwGeDvA07K7wvWcx8r7BjFcakhudTJmMUmtJem2scfVtnpTyGyULaywGRXtS0vG6WRo
I0ggknmZqh31OgSxA0IYl3OhECoHwtP9S2sSvVbJMwejVy0cEdax7JPkwx7n2ybWtn9FBGpi/Y2N
4ggDJ99IasFNTmLKII8wJnE25bjo7Ex9T/gFihCYBR2c9ZZhxKg4ev2aSkYIRxZ0A48IuguMPJeh
6Hez4G63RNJpwjS+apDdlo1m7BNPxum5RHMp+yimW2XJugnPmaUd1JJVXyiMA4q8nZ3rj+rdEiZH
Mkc+VFcBufz0WavzwVPIlVGiTnxXEr/yOj1VXDWtYDY5ekuSp1RXNDxxewAZ/3q7t6o1pAhiohlY
u4yLJwJTvuZ5yRjsekQtUo8vo8CaK8Zip1Q2bNhE0pJdzwmLrj4pKFk4VsrOpgoVOWLfApxzZR+d
2MZbm6RABI6dFJ2E8kZ/PGX7Blwq08WEpozIVF8YeWVgdmMGKGUkk7yGFA0vfQQpWn8cC5EvsFWR
Yu425WkTN69FuT3pz6bLbFesAg2ya8+OYPuOkm8S9mgQaxpfamYYEMQcZ2ssj5sO4s7OirRe6Ko3
C7dBqGNZWH8nWXtNgOJ6Ykr3yQlxwAQfjdb1BULxjvWCqcvWWr2pOn0s9NG1OVJ9xTPXjiBzX+GU
7vMwkv0HvP+czDa2iiLPkV51TSGyRAucmCoRqGbrFBkLzH9pLMYqkQ2IYmN8BAaETKNAudaWTbcQ
GjXAHDuwCqKDxPf//bW76BPKBi41HUmmBIFNpxHlcDiyZlT/Nf75Lbz6sx1aDYpTe3P+7955n5yW
9syEbAiy0uDAp6dWXgt1QCsPgzP/mH75yGso8WjF6FleabjXKsTsYsRKUy5ukpkNz39z+4v+ck/s
IGort8YaeXsIp78rTFQXyFNab3cutmybWZSpUraE9xmx1SsqULqV2uZAHMeogcwwc0L/gQOI6LpG
AXlYBUVsF+mFyBAIOe/nTUqBcQ0DBc83wy59yRj9NT9tC+kQvj0Sm+mk4x/J0o8DzXURl4MLxfsp
hY86JMjToChVWUFDDDcXoqVt8/kzB6XEn9AnVKnQ1pg0JvDb54d3Nv3Mu+doAHvSuxlsZ9wIxW+f
wSzepqhGqaqT9UKxi0ItE/mXrIyIUTYDFQSxerBMxdLQqp0DN3C63fyt/wonZ5hYQkonkH7YHlAF
vmaQ6UOwHk/kI6kybyrPL1TScGtWq2Myo/b3pJ3LIjw2kpD2eG/nDySLCDhZcaKd9cMzlivCtjTM
Y9FR2iME96KpDryYYoWEC9OEfZQ4fxpblpFyy8UIjnZQZUyWnDDzcymhxAgLs29MzIQcAf+m1MhY
uFmFUdmjwCigrj5RZ1jx5p1YinoYRAg/bxx6fFy9TN2jBYYF2tDA5JZn9EMLDpnHIKn0JaRamRGy
YuvQofBE3SiIk5OWBYtzSZ/WwcU9O88WxEHnFtGV8MgDQV7HivbZSyh8Aj0oS8ZU1PKUkpJC1gUA
QIGPhRgDLrrcLJykvb4A3w+gUS6Y056Y0maybq1IdvSBgDiqutwJWZ9j4c9YLI22JcmmBx6nV5UA
Z7YGIBxNchdRC1l5lePUNiV0ggEqd606Y8e+hzZkl63Xg4VVDtLCQbf94RtYxz4+ueTAr/KeEH0n
ehnun5k9iCv1Z4NV79Zte9bOI6LaZ/S6CaQ0wuDfe0LIH+K0q3yzbm760Or59a0EX7zjKmN/qmGT
eqXlE1vEzfFqHiFgCfHtI8nR5eKp9EQN4u+yFqG4Pqzt0wvnQlnwoqS5SnqpWZESstsBVf1mdg4a
GpdSXcjUMieHr6lFGFWy9HrL/n+JBRpZD41mRGElOhw38ExLuogHqdC3rkO+OcnIV8NSzFAoINFv
xTqE48X4ik75bVCsjloePDUGzSWKIIMl6P3zA/7DIUTpZ0UXnczndrOYYXC/YnEJ0WsYJIgD4tCL
2tDAhJFBzIqOF+4r/wN1CvG9hedokKY/7kVIlDBHfHVoXDDkKtNFraM8AOlwKXc+HP+QmWUZT8d0
9VeRdaWLEULYFUocSeBCJhlXBFUxkFcdrLnTuXRZj8NVh8q5mZ/X101Yn+j4ALjPpQLhUwPyR72p
HWVt79Z8s9PyMLXlg7Ps8S+x7Db5OUleFyYo0Vfomp3KKVfKawbK0clOA+OQWZYYgbRXWlcA4nSx
ocR1esRpaV+2ip8dnTojHK464sJ7xp0QnhsYlp75xuUba9ySW84/w6BbeqQOLIaEoQIDi15X64qJ
rvuZMVtfeX/vSCQqUFvAK76EcETu/PUPBWLIF5dw7uozL/JXgExbAH2zCC2Hh0jfYknXtnzFE/xP
3gKntt7OQPkdPu/2BZtFfZQtpDs5jnJyx1R3XclTBKC1bFksqnqWIMGIwecGhOLHeAiBiC9quArb
KYaH9DVWlhqwnbS9Jg9L50RmTZMcW5rvPq9p5atlGiLFdHceufhD4Qv4LeulPGNF0KECyhG/HiwE
Oh0wyWFCnRVJa8uM3Z68QV2cNJXZUv0avXaiKxgNkKlW3/18/PXA3BhTvvczFPsZk9TTmm20E94x
wMTCZeemo9jGpXUp8MiICZinCGjtN0ro/0HLvm3Ew7NWDUcFpb/mYDYZ6WSW6nq3GPyAyo8ZKa+/
fWrhLf8xIziC5FnhKaYncvmLkqn32YVj19twu6y5wwo9TZEaspkOn7UXZhVvzP3azj3UWiQNcZB2
vexi/Onp+MQXJVIJBFrLLF7qCQO15GYvR03xgibJWVxpZGcMUqm04ZJvS4W1GmUoI9pCgeCe+LgU
TV3MZ+QNWsw0NaSdhW8vtKBATo1m3g52CSHSCejf1WN5bC5X9sD6AVutXaySSRk2SWzF1dCELuH9
nqzpK+SE6EHDSK5X9N3woX3liCzOBu05IgCYoHM9sHuhhwcQ5GFYcOt6AGa1b2lTMqUa8GDM23hn
kyFO/PpIvUOCw1/DDCRvj4h6VgCDCbRQV70Lf5oDuS6DxDvv69Wz81zZq1eRNAfeGiuzqM+roumI
metAj0uVl2nPAuW7rAyB4nbU08FP5yMye7D/v4hvnHwaoZZPbgIhXadAGPOdK64FmXzwBkcWRgxG
JGe61YsVV2DlX/lGJVaZKGn/ZOD1ULIl49T4ArzUSt80hSjvQVRWd4s8hkbeSrksDqnlMvfHH1lS
JfkDhaRsQszo3mP8UBZxVuBSURaEyic7jewsjt9yLFYX3DsL8pUQA1HZlvwl9r4xGZ+KGJb24smI
kc1AKSyjU8/fnulebB11zGCgFhdF75fqsE2nTJCJsWZT+KvrtV/cMYYdjnxdPf2s0MJXtAfKe46g
yB+Tk9PztDYD38gLeurPRuzkPGkEgu+LzEInLCCGf7FovgkHZQfl5SOcaowiNRKxACRmz2v9CqIN
MHfNrKLAMZ7Lvu4kYxx+7d2L9IfxQkAqjaCLirCA1bXamIVDoAf/13UsX/dxDbK0nkUUXqHl+DAF
nkOdwwMeE+sGcyPSp9tYebmcGNJPIl0C43Ornq8LwildHdJB+WOp+latvW56q0DXS2E/b19jyO9R
HtHfDkln9cpW5GDN09ssSROH2WDuEfJ5OpnjoLp427oXTeq/kvTtrgKywC2VSDOB+qTA2mn1xh+8
utonC9fLLEFHV2keV8Q4tKYBPn40INm5cVKpDU9cbFOMhcLcZKSzdrayMj6BedjFnPS1k2oiDhF4
PravLzoPOcfvvKuvRNXxDd9CABjbP4KNoaoR5D8bJvtqXjJRsE0Ci6P9+v0Elu0d3VZDSq2vVrXJ
twc8dvHoqPQJgfKMH0BRwo5z24Eqm6jsrPre2hSRGc8SXhKL824BImSvMqte1939GzMbOVz30wWz
0gS/nU4C6rFXDlS77lTh+hNPDK08sn6A5HlpS4OU91ijlRtSzgLuJa8zN8dpdZcN2GY0hCtCJVwr
rp6swNroEQ5NKv5r8HsAUxahEhEDIHDql0PwfCRCJ9ZEGTrzle4k0NfKeNiEppKjDgYAYJxMcabW
DBcmKDfzHGUZ9XmJkD3F7D6qzXV9cTfmCn8QIGYF4YDbZSeoxu+Zsu/v/nV595UN6wE+ovu+Fnqy
IJJlT9YuQ19TV3be92uQmFbqf98WSi0pOfT90b4Xprol66hh2spTBTncDjTDGukR+2TzD1L8/6VQ
pC5XR50tGlAV+zJ98hXoBg7Vcroe11m8Ifh30isVm564IqeGcrrrShE26R5uMtdCffxS2pjxR0sb
tIGELngIkC2pLpliIqKgixgvwoWshV7Ckf4i55fycd1NGp8f6jiICsLTjoCw3SCR6WJWGet8ZeuS
NViWAyknCN+5lvOX8kGyCT2dHAKeDd4d4XyC16+ianMv1JFAGmFqw/slLdghvdk704brvTKpoaFq
aOEJuRIxFB+dBNplouOwreNUBrA2OyRr+ibOS9OoLltmFyPPAa26+UOXeL5Oro142eQ2f8cQrSZ/
Tll1X1DRfrrYOQ1G4VIOo9m4XmQUGjSCVGzelt5xMSLbCoaPK+nbAFkkazRr9Ep/ApXpbi/FjLe8
rIiVZjnf9aLKGmwVezOmXp0M3mnJQVuelkewCdv7qUjXeKi8/T1QV3T57iV/lFahuZvkYFR5g1EH
JlkEFBMRj4RekvHzNMUwCnZ1DThMJloMe+4TOSU2ZJQ68vOOHkhIzWTaQgvsqLkOGrmVgvQJxIRK
XfOJ6xWd5FxWmHXgy6O7i/8eEoZMHBdUCBtTjQgIM8DPyezAL6GR6FyHT6vVBVjxMBGKrhw8/fw4
JDyF7sGht7VwX6gPbbD2X501G1+niriVjAzP9EjMU1v3r8DfMWYnZpXeLBh/+su2sATvb92IkxDh
qsMG8JMd98+/pLoR71sCJ8nspls2v3O7PLhmlhv7gm1tXTeS0UXkJZyDh9NJG1yP7WGObJssu9bR
tAXUhMzKrIKVpdXWSwH7ViS+pVgvrRr3PkM65m/DfF7KA6vUHKiRa+Xrls3dEsPPt+VtDaVLZB+d
uY1iVQ7VZSYlup0GMDqvzH2dNqvkbFa6q6icl5ag1XoCEbzXi3AbMicX34p/LS5Y+UoMYii8fBkj
adLwxxuQ/zMRX15D9JeR9A7hkdnAljWQIYrxNzhJUajVLBhVNw/ZmEHISs6g0UfztQDyz7pRkrgU
reWG0+4erio86fryjEHVjmhssn186sqVIltCGRBHHq+3+I7yLnIPJKiJPrcIaGJAbwfxadh5Ko/5
BM/8GtUaMOcdMDPpvYtlkXz/EQm8ng2OxypzZQa83c1Y6SBsR+b1bNIc+IDncseyNQ4ndXuemZJA
lrbckgxfa2GNzbaHiHcAsdJ6BMg/rZcxxseTVJeJDoqB4m067oAKxDnSUj4EdkxA4qXPv+Zsh4cg
Fc9GcaZobfd1G/MAdpp2rcpiN2y1FrcMuH1Pjj62nIu8TFg5Wridmo7KD7tFmOOxJf8h5n8euXKz
OcPoUAzlBoX9W5qIOsBAyHpjC1WvNI7JRmI4jKdgX1eGgyZkY5FhxrDanmTX7NGZLb01t5lEV+q6
0XxTkuc2wfIaNmb6GQYzx2+1DC+PkG+Kf2E0Y2U108Xm+zw59R5d4FyIzLY0ZkJNBoGPr4c2jkAv
EMvyVonUrugBD1xmAZVEua0TmiRlmFvkYtomTh932Y6WIgcrq2WJk7QoMz/ul69ce9Hqk5T6TKHw
ZO6y4H3H0PQXF5xdsKtzzPOyEJsvZ3HB2e37e6IsLB/rw+7ucbcyvPQI3/uwfq8rVL9+FxHELyYu
h8zs7iXi6GV78WDS/5/eAfGZdPePhPqBp29vE2mfIYSqZLJCf3ET+WSmecQNflbosV8Ni9WKCn0e
n9daDp01Zuux1qVcJSO/KjPc9KT06BY5KbffcVUsefHhw6mbjRYTseAS0MA7gOmdKOVMk8lWRgXZ
2VCuD1DmgPKixpjgDlndWxptXCS+p/hKgOYTxPrNMKfQxW9ehWQqrwCbiVhSgAHfzp66QocAXh5j
zw8lu/V747ytWuqY1pvWrs9ecq+mpf2v5fxlX+ZYrGhgbi+1loR0pXchL/EPnj1ZmpC/2jHlpNX0
E3DSgd/L9ofFc9peUbdOy2FiWyrq8mKfl8Ez3UOOIPLTD9z8WcDfhjtL6QxBhcwbSN90RqBtOifu
dxA5+lk0NwFADM6+tM4o4bPCnp6yIVFlldBwB+7Sbc2IGqT8LFbVL7XgEtK4Fe2/DIV1ksxvTNU2
vAzoq3s0Xz9UUAE+vDJ76OhbEeDOBBEYuDK86fYFP9C/Mrel/Wv98ob07vViqiGDKIiNX2+1QaYV
DnhwURq9GowApF0Fl1JopC3XCfkwRpuTUGgIt3NXqnb3atd7yjiyjVr2FZb3z4MLBLC7Vk6D2xov
7DuYRKUKBSLmIaZNs7hNPT9oGh/xri8NYPkOZC4EF9tbgpNyhvH6sxLYo3tQNFrthnjuOnCP3ZK4
9BLv6aOBlT6FDtZp+jgdnwdfZNQKJV/VFf5mjNM5NdWgRzXrvo7FOnVrzwm7BnMQ4MfxUCOJnzVK
eHvRqTht1KrbFadY+S6Fuo1Mgb7Y3cjby9ojwyBTbth/zQ2S8q0H9Ceo+knD+WqcrROluZnb0ag0
mcFZta0akhUi4bmRRAvbOj2XrW9E9dV7KKzMVwNzItlTwmCu7ZuTC2mnI5IpmGCOc9EKFcxlaMrv
oqix6lT6JMFayFs39HTGAQGVPrg0QvFqm3Tr8lSWCh1xHSPAgmjowTBl6wrXSi05KJWY460m1geW
6mBGeR2rz1HtFQXtDSahVMGyPO/t85vcq6EdNa7M6WqdzJUK/snxQ8/o/ihtBzEX0axDD5Kicn6B
/iC1nK0Ynuc3TVOl9n0zL3czy3BlbwZnXYofqBJedP0LGQu0svSVtYofg+HUaBN4AR8LV84aO6QM
OAMzygl6tHT1iT8pFUdDzF90+6fdSv/FTJ/TA9XQpHfVGfhF1JoFiWU59m7/ByZDCbBihDugQIK1
88kjz4tHdLpWJE5daednfDkUvcF74t6BH5BTCX70UbaOeuRbuSqhIhqmeu8KAPUnxJiQQHHaEDrL
+Jhbf6PW7wUNawD5lIspo/pqhwE7DcD0PtVSO9Ygz3UrxPQuErJwvDtscF6kYRm2IKHXn604mjbs
bhItbw45W1SScKtN/xxgb/biJYjwmpXIZo/lSUmeyoyxYCgQQpmWZfTxPTVd6yNEwQELgJ5VLBgM
LJ9TwAwan+6K535xiRNmefGcsdB1oJ+8PMDL5YQOo8NOLYWL/oaZLCXN9KInFNlr5yT58uDqN3Tq
2e5FfnXOSsClxOnp2iNnpYCO7tJKXe8wVXcTi+JUML3RH/6VWn4LKM20qp8qS5EwXT22VdNSMPMr
aJRCJ1EYbq4UTFbkyYHQkt9wqrPF0FQ3a4K+6oVxFgSU0+Ynp8XVmRqNfOUmVkLia/6yFtRfytFz
N8TC73L/a9CA7gJpNou0rTr9AhkDVnxrxORemu4c1/cbtN4IKGu4V8Gzt7HORvZCE3JE2pBFYcz4
8cjy2g9x2xWNJ3EKh6I0qxRAsrWlxuW8zq8QLPeVlBSPDN7eDBZLDJXSIXTjOtDO04ARa750sHqd
/8r/6w0FVWM5637+q4np8jBCA+6OUKeWUXn1KOKRI3OXNMuYCgxt4D1FSaH0uien8BN33SvTjPhT
mkuDMhRQVatqakZA2TkCglCQAXB2kVN2MX2lL6HaA7BPlTs5IYIEkdH3okRjXo7SzIS77tljMDv2
RNsC+HenkRZTY3rHIBthtXN7QX/ljBYlfbnJ9zkGv/E7imRMbOPdtRvbEIz7Rtq+M2d6ZO46b3ep
TX0IosJThCG9y3cX5tD9VRCe6iYsB3kLGU8Y3Y5W2U9nBmsyp9XVZg58GyLd61kaTbZz/4vxNXhb
GSyYygu59BTosnVRAdDaoy9eUdkpT4ng2Q/Nt1+virYYP8Q7qxWfuO9cYXn32Q7yGniZDL8KO0P3
XW29B4xTq897L4UsqYzBes3oI7JGwdWWv5xO/54rEJQQjwEzd3NxNORO3wlmq1gXmYrNGZ2OSkfU
3esXUPPVyCWBpICrUnvcknAP7d7DmyeyT5MBJnkNQzrKw0fm3qA9aXfmw0sVdsv4EJSiv7dDCLCR
SlhX4bg6Huuh26dInCHZvXUJsvIdMtLZUp+Rh2A+wr2KMNXp9SwI7GUlz0oAKm296vgLPZZdUIHS
7xOP6zXrNhoBFbhv6QZQ0v3hLQo4wgQzQXeQKxyZ5fyQ4h48Qqe3elqMu/ROB6Q3BnXvSVQ90cuD
3OVI6QNKAkzxON+5gtpOpcp+gRZn/TdCMlnlRNXBS6agbLpwIURT75aAjf9tyIb9UfrBCJeCTYDF
0HocFJM8XSUMqelwaufPJAtoGrKWeFAzQDGDj24wd/t58mEYTHji6S67p9u3G96sDBhAH2kv3Ek/
T+Phwa1zyU4whpvxymjvT5lSFf2bppQ0Wky2LMfcV2NE1ICkUkuii1aqMGzb8C7hVSmGQ0Q9wsqv
osRN70KWGPyIzUewH0i54j+X9uMlMZ38h/j8izyuQQl62tezu4mSjT6j8NAYage2PXK445cpmCe8
oRKvX795Pk7V5n8U8YN5ItPQJ+CriYxXuF59fwFRKUcIUW4eS5q3bzv4lOLH21A+/bho0ExuE6pR
4cIbNyFK7GgeCDzJThHj8QvL+SkWSVZ6PahIrptKNSj/FUFH4wbC8hLCrLnCGIUCP1nJuJDgPjZp
upGjnEgF34GQL0LNttMF3hM4VaXxLKLnA/o+hUVSJIiwLp2JXhf4xfXe8RmdX4v97++NuQck65tm
SoC4YGFUx8jmPIIShcX95BTMZt547yxPj2l+Mr+ovQX/P4bLE4hine5qjEPpyNXMDhhCEuAyfCNE
lmlgyc7TirUQQHjZwMVQ9cPX5BtHIF+KXpsAZW06nY1LFL2JfVMBsz3V7wGED8Z+laiintwt+Qjl
MShUVy6TWqJBmS2xY/bYdNurTX80m3cq+9OrHva5NERWVqTam8aypEZl6lXgCqSEKGO82Z36FzZJ
AjFpy1EH5ZuSWwLddhI4SuRQSVDB/RwW7K1n8kgC8RIZTSfLUHQFGdMrT+8Xhe3AIELa9yj432B2
xVtSxnrdBajV0rKdT51bZbaVOUtsSfQusd0uiqsa3Bl12noLdI3cqkBxJ93ZhXUqdQF5Llul1fEu
sKIHpmSXzBIRKy/SqdW3+LdmD3n3nJxDWUPhnyg++PrTYf7WiV2Bo61cfhEJn/A1aP3+B2zmzuQR
ZbOU1gwNoTkW3IefUgdMYbHtYfpsDo0i1+EL00UnOzgZhZQWUkZ/hvJO8scbqm5cKl0Cr5D4izo0
2FVAJ6xR8qmD8yxJBjylyediy8kE938JWqF3dT+rLQYT+PVvu3hap+vhq3Z8ZcyknAniryFCuoIm
DcmUY7Q3y6gFLurM7pHptEDPPzUt6hpOnNYJqT8toxLxayZyud85UeOg9p4i7ZkMDfdi5lRmYeja
bntek9ERSgbKUKC7mk8AOVlpdDtHcHYljL+fgMazufVaqzk9IxUoR/MiJdc+8JLjeXzFYyy7w5Gl
2Zg9HvgnJOjKmahwDTIZgrUW0pDy6h+nfdyf0KiHfLJ0XKWYl/9nhhSwNyL8Xw+44zO0t2tdJPvr
yqXZeN3MXHgCC8QFC/HMJuE8KnledDLjXpxDAyGLDyrLZ16l3RYpNvXbaQzSaunFEJqU/gpdqL47
97NAtrvdqGAv0GrBuqJK9nsvdbFI2TRNI/iW6xRdqSsxZ7bDisvSDXIR8hJpDvAiDgEnhJHsbYii
O8AAvIgR64JU+XOfNXc9Z9wYJ2Hm1maUPD9mdZVsb/9L3Gbuvwqj8pmV07Qy+ZX23dIbKgFxT17F
qoi0cI0Y/kEMK1AkTOyJau2vkd8d0b8ATHnHkTlwrGnGMA6ObAZzxXYj2z2RzXIPVTAyxXyNMWIT
WUkEB1ssC8ImDayB+f1WJ69Ry2Hof+v9h+kx3a3OgZyFkzEgNWJpSQ8cjMdMZoFZzY8Q96f51hxE
rP54A3AF2AsvGWhCdfWqZLIW4y05Yeob3nxurkYTCIj2lr8/4dt4wY1nuoRIxHglRli/byAYko6E
yM5mvS5gJGmRPmX+AA77DkHAZMEMEVljqDNKJQL7G7MnYdAMB+BM08S/fbORHEy+najKHwPVx2Jn
GU1VDZmAuG82z/87kGYfFAkmwYn6b2/0KhKfq39kPMgPm6LvGst/lzsRBT6gyj684Zg/5hQA5PfZ
C5EpySK/Vzk3sDffLdgOxfmVMsn6IMa38PensaD/Ma2SiiCzGLDJUPliz+5RxSJ8xW+KEvFHkuRL
W+TudUnH+EV9l0n9a8zBZc2eiHCGiGmt60T9j+8Ah0FKtV0zTrptbQ4NlV3ms7YKMfe5EiKjyRXo
JTfJxGwbGkKIvwz6WYdpWNSieStBBgj/yUsz67z4oQmfQTvkNZNRsjgCtcswsVmLjc+2gh7i7bX4
c2abuLLpRW66cOHWWkAvk2Nt7dHflTNSCNvRA2CaSV8mq1ZRz7adRvxh3DwTXmYK6ys/UDIjY+ZF
fEUWwcXgNNhNNnlvELKWbDpA8P+1X/Mm41MgOAACfDb2tWsZL4bWJvBFwqz7mO50uh0DF94ZErPY
iHy3ttsapZKyLClef7WlOH7nJAV4O8YHPvF8YPoy8ZP4/MPpek49bnFwiGNe71GjGgNLSV3Vi+gF
6so4HPz4DEeUlgXYKC1nvF3HUU4c3JSkjF/Qc0LEw3hvMR9wIoSUEjlXQ0LAuJS5ZUd2Srh9thnK
ZuGPKA6Emfg7r/jkvABjKw0Jl8H2iurjSemZM+tdpcwnNn1wQO6YKcF6jXZLviga9360yzpovGFF
YWoq4/EhZAB0B+7zGXfoNeFcFNYQTaxSbsmTDy39fGOmRNDjKpt9PsVQgw84VuR/cHL7y4x7xoY2
3hY1/R1GCpITAcS6gddi1/dol1+y3z/fgIZjSnvwRJYYjTukgaNHmvWN4JkuwjwwvRZgcxMJpfJz
i2WJ5oONbrNLjD3/MF1fvRcn+fqGirzD0F4eu/pMdu1M4Wn2hE826158pP63m5EQsNadoZft2vGd
DtAQ2pWmX19PcYmwS3RyXbEj/IkOJrULO+6G1tCYzlqiobmkJQ6MfheiBsNd5SepKz4ep++jX+VS
w87QMxVNH5lUrn7BB4hKpewHdUkicKD9A244p8gC3RryfVt2gt5g91inlpWgCeCxYyis4cxx5LPX
ReBR4Mb2tVaP9fIQL/dFXaoOz77+fo+d2gQcAZ+bSFQzjjNDYu25zDxGWBc56667DvbSkBU+ftTT
wop63LEoeYPnUXblxINqUsxhj8oDR1Qk/7RD76+5pFxnNAxS793+kGK84c4AddGiFJazl1YQgBxb
yfK8lFeqwo/ohD6RCaG2S7Jp9by4oY3X1BHA9elU7tv/La63fP2OeeFBvO92jHmHgm72IOch8V/c
D71D6vXd5CjyL22HQrCW8wScnZKZh6nvNoVRbpuzP1Ab/aNhch2YKtWcjE31KWL72Zhvl07NUVmI
ZQMFJ3Mm204DSI+P1+6abqNEiT8stnQjL5wniIxOuvS4QVMqVw2hg20HqBGB10XllERQ//2dyMNu
Qny3Kjs3eui7Ec+DSj3dpdp5Gj7PmW8WtO2HC103GMv30sJPcKGdIVeOudmHd6NqiJcOMBV9Vy1E
UD6lLG21XlMPCBPDnmVTONZBUepcjM+M3KFxp+QFneObHwpM1SIEX58azCM6kcyR50AsU+R8M5sK
4fll7XD7eT1Lc6O9v5efphMME3Ogg5+YGUlAhVoTnVscsnyO0/OHtpgHNVTvfoY0y1apTpR31N4A
2y32+OFsGbfez8UGANgUs20ODBXjhirZX6s1x37QW0U4K9Jhx6kvQjKAmdLY7jGSNVkurACVu/U7
lmQyyTwt+aU1xtlgejWuIB7mmeMLbg1rESN2Ou3t6ffcKWMFJYa+SxX848vU49qKvwMp5ocqut2B
QQFK0EI+KmvLkXQr9zFEyqkxpTsT0YsDA8l87ZiBzHb8phODmZ/VFClKo4/xn1qdoU/MHq8NP26r
E+xFjfOdfhvdfLMp0yfuFHCEC8Gzw3PR3f6u52BzWfok70XZRBWFlboDuazXF+c7u36e6KniGX7b
GcUarYhuYPBREnN785DbwzNgOaWIO6BACjwsSXPa7nXwFEnhgoeBVsAMvv/col21i7zKDV5GTCtv
I9QV0ZUrwCd9ISy62pyuqCqEpFH+4AzdTT7et6q34Y+KB1LHEG9i+xbNlap66Yv0FBRDUt9MqxkJ
M5ivFTXy+aquCEghxf+I1pxGhZQHf/2ZOMJOHmKIy3Fwd/1pT1gbZN0th8bpv7bWacev8TObabGJ
4ewCFt8h+FdALfi4h145+Q6hF5F4fRXZ7HpSQXWj699MLkpTSpjxdrRr6Z+GAu6YuVyyOLhnaPpn
o/ITgH8IWzGO0dnTSVszjB1Ua4GraI3dkxfgzWuyHxUu9n5/WFpVfsHGd5r8AKQ5zAMGl2DMFU7N
WvvmIQZP7hKeCxx8aIBszNjEAuCjKybyddyyaTpawEqi4JOta55ukoEvNEMXy4xvaT6KOI6dvywV
MJYR3bPsl+CSpf8zUvV7zLfqpGAi5yGUz+if9M6M/Ym7iLbTCMeUAZvqv7yMzhsbcMAZSCs+wxV7
2Xn5fTe0RbEOC5GQPOWL1V2/ZoDPcgZEV7pOJlgIpA5uEWRgBaJWOx7pBqc8813dEHToqWah+03N
e1oltR75IzbaF6rXm5Eop5S+B7CTx0uADhhjYIldamTPo2akr5EgkhBCV74xntFH16gC3/Laqylc
Ietx5Ha9KpyLfc/Dst4uz4wDbU0qR0G/BglCOBOXEeqoYP5Bj3Cl5ivulvUniYkbaJfLmiMwb3lj
OMjci9nj73ApH97f4AJ5kmHc7TInEb2e1zYI5O/0zsIP2Zkk2wzeUkNBzJty41TleZHYQ+GHZY0D
CqwrPOBa9oLankdklWkgjjgSgyTbAx3pEXBaYuL9mdaJN+rwVC34WOTHRT09CrOeawtB4tluFC0b
KsLPKpj1fDc1HcDjChAObBcxtuRca8WmeF1AJd8pD1VTLn+D3EejQ00HOWFWsKqGcfW5Q9iUzBnj
BVYUrRESIWzfQ40n1OtES56pqLODoscD4OhJl7MMsGAXlDyYrcjFRiC75/Vcv8cGqmHNO8KKGSs5
VlHQM1K2S1P+LoNnH7Rq90I6n2ly1L11pIedQcGOVVGdNHyoVMhZf3f3BLX4U/YWzBH0Grey5mOA
9OGAd7XCSC0+Ijx8pja90qpEUgkeVl6nfU2HqHHhsKwbI974jIyT+EarQ7YkuUp+/2Vv2zJLjNS5
OBEDegT86t42V2qvmg/l0IOfiMylLEYkNb4I6iTIxrmu/T8Pw3FTABCiPdTdG4JmsDmbiBZs+CR1
Qb4dS+rFSYLi5FIjg2GLZfrJ/g7rNsbsa7U9lM5+1/7v542S9pcC1dGP9wKdpGCs/uQY7xCa4KYl
B2rl0dYe2r8KJtOOtCHiR+BBzwdzW3dNb46xBTY9S5ghJGPP199t/A6A3I2ScrkLrihnoqUV0Ms2
8NW427JPM2KlQIZQTb6bNhMHNSLIVCTl4ySY+Lpy1Yk7t+1jd37r4xwtAYW1af3ZCzGSQ6AACcpE
zZvnbOemJk3rk1wfubUyFrv2HTN7CQvfK7eXd6ohmRf6ZfyIlnuN4sN/FkRicPYbovhhssbI1uJY
m9d02PLQQMU9W8UsLnUJogiIaz47Vi7PG16iNILcrvM+qqmkd1xFXpK8XGMPWXycziLTPdtCqc8o
9PlwpdCqA99HUwNXr0AcWvP2kL8Yg7tR56o/eOTdo0DNj2xW+SgH+T7MI/vwZfTmbGf4KJJjVQGU
8yeBPjf5kSrWqTbH+rCNYlIL+2dFVP/agcNwgqJdSx49FgEM7rrFPhY+3q7O0KmKnRqoyrVb/e0F
ksGWkJIwjBnyJA4Mq01YOWW5wKwJISk6wGMCZ/qkiluBuA1ya/KYM/869lTsWvs6VSq4Fw4IZ+Z7
bz110SxZik18MGzJbIfJkKd62CbqW/yWZn2VLGAI5tBvn/YUQ38jX1xYWUTZUXUk3fq7rfmDwaKj
vfo5ik4M3ZB7CiazQtW1vbSq5Od/xcbe2TCkTCyoBQrURruj1mAGIRhZ/dJOkenqid8grtJZ3DCR
RpPiegFG3DcfXFwHoc6/vvZzKOk+rbgacqbYFtYBjippvdGO+Jfy+v/Ta30ZgZmbavbvTc7v5cb4
+ptVcHUR5aQX77D+8njacuIn9o+1HtoD8v9Mjpw1ijZRi1jN7usfGtiHsb1ouDBf0Oqzan/pPM0A
cJExoYlI0Du8h/f2TcOTQA6++gTGQzLen+k0+m1XalJQKd5LCLkL+M7uaecmrbiW3iwe7+k1qN0R
1IQbhvl9zu3bVbDpNZKP9TgjQvb1HAKUfFI6IS93G5e2syuYFiCNud/wcV7KPuwuudvbfe9C1lHa
0Cs8I57vViyTZvdGoPTFVsEh6YgLuMH5lhHpZNCOSqLgYrR7XTNpzWMBggGCoE9ePb7DtZlals1n
Dh0Gze+myNtbam30hPfbDVKa1gV3A5riysS2N7CL0kq7W23maifl2MXl17ZHMylwPl7PFVd8s4gF
l4ukhZTm/B66OaYVNlMqoyzGgoh3piZaFfZYLVYsMz6V/UIy1kL6xElyZB3+0l4LnDm0UcT3ByLf
HSUQj/2+f/Z9rfpiXOUqqrtCIc3Hv2PMkwPjXJoIjBAxV+8B6jL0DckrJn6mND8dK4IK7OuJPLYm
cGBXtXuEPZ289YWVb9JKWyIRUeUsdQEEKhlDZHF72XbuN3J1S3PPha1zcTTAqdItjONaj9bSF9O1
c2OxIPxdeW8KxEeOADyq6ixq5aOg2TeU1xTdsZ/Cq0TkD/fjk3cVWjkdeVEDFIzgdK52eDMpH3AF
0l57LQ9O2S4oBXYbJXLqOHwQHOmkeQqnXukd809OvUjVnXQ9mE1hRDXPHWWL8ENn3rdKGxhQ0Ayy
IqKiojLOD+pc3wUOKQ6JtozuRZVThxcPOs3mJTW3vV2V5PJMZzfEpz0xN3hAquW+Q3sfhnZLzrOR
32ct33OCqndewgzrBF4Fgi0lgJz2ctvTqJfxR0z7XQT4ya5EgJMTAP7ngnWRrq6gkhIGrKh86UWw
j6XdwY0I1gOq9OArXeKpYRRcBTXKnxLTqcX827j4KOTD2FvmQ89UZGlJiwGRLj+/trUBrLHpm1z1
5hAFKjeYLW7kdjLj55h381VvjeIO8qcC1pdQHGOym92ymZj0qow6FaNKVOEHOCOGITDo2B/TnGpy
ZXZMDKVdBZJ5tf6Yc+mVMptuZLJlkzFj5R/Trhg+CqJAw6D7n9y0apH0wQgRu4aRyNHzUnKPZmAC
adr6zXmXy9FqzgkJTQwZqbiQP/zNLr/KhYJtaI/3HTfAHVssMNL5PMUyRvqrELLuyBpG3YNpwkDI
6fXnJtiHgDLVh1fX4vFORpP282owWhIcYNCSzIL/8HAw+qGLITxeM75wVKHDrTt2zNLIvcLkk9H/
HgeM09UyKZ6DDUzq6T18lZhstzQJJgoGTfUOOOCgZnARIuDgghmFS9loToN/qPumwVGufxudExsB
qQxoTGuQBhLfk92n/Ts6NvDXX33SFlb2D744NMp5NYICkb8LfSsy+3CKVDVb9T94li0SLBnvACms
r8MosOo9+Syx3jvq9RqoGsOVOm8QYSgyFwy61dUZ4boaKqHddBkr1lDGd4tH+4rsQ16Og19Y2U19
ooCn25lIvBd5FN6HW1B694Q4HYbIpo9eUhj9c1r+r7uDjxXv2m7vLtKq4ekEcthkf/bxGQT4tm/g
T9nOQw0VA/M1WJdGWyjIVAo37RAhD91fBzsflha9bnVHGtNAQrrJqCanmMvKaIAFr3RoanmMSvRH
dsqy7j4fk2vZ3la7HKaoOxyQOH/mY7+Fvu+/DQLTCyGVXgbtQ40lf8dXIrp1I1VtfVy0D7dtkgUs
4ymBF484L0TX7nVk27FJWodeOAnvHhSHr7nDSYNSMY9VRtwK6zUrejjcC3YDqUyquF0gkO8hzde0
RntrJVs/AHocge3fh+V0JBjLuGHOK6fOY26Ls7qiujrk1gUGT1zztrMtArfgm5y1Xi+bTCRfS5ui
rKdyct4wqKBbsT6MCeYHUXC5s3baS+Hpxq/FoWMd8B8xG2tecnMJZqfJdqMcriR4z0YODJ9yZyAL
6PumQs5bj3/MLWuovUU44EUIvrFjtH78T5OFgfRLsfw9H1ap/omdgg0V3d1sV+3DaPjInBYt4qHD
hW+rivMAO3lHTLbt6thok4D+FLoIUkuPb5idOp33QyiOI0NyK1hBreHjcVyippdADjkPXiXQoeky
gHYNDjS0HoWPVekN3+ByUDA6Vr+1DmPZM7sFYzHNmbnRWRKfjI2S6ljXwY29fStznaEguIx+89YC
8/GeFP9v9ILLYCKc97ZOkVBTDBA6qUX8J9bwUECy0nOX87YSYc6VJwTHmp1itfh7EyWpsOzWHzQr
agQ37J+2mQq7g8AHZbAAt0B/oEEzSL1VO05Yx3T6MXC6KCcL4M89ZMPlK3nQJM4bnEBsgAynlOet
8p0PfmtKfF+0HRBz9JNlLdGpSHOraVXreaydABI8b9OJ5BAn6L2eIBiOc+7xqdtaxs/Smb6Ke4E2
kAxq77pKSAcWrkxp6QRouDFqRX5BwbUK+G3aSMmcylgHxEIie0IUd/3g7HCsCnhx3EHYrtnCmN+L
Pi2pLO56lkMsfwY/I1beZr/Zvd2kVgx/pmUYELDtoiudBfVYkCcovG0JQHnjinlJerrqs+rSXL1F
sUcjKPpTn1ooYoGI09FzVrrGpnsdqcTugxdSI36QdSigFACCHJJiX+JNj/TIxaSqUY5rsksE04pY
hXclwVoLeT4bdVn8ZP+bOsyeAoFYfvIIB7gucdUZOcfiGHSj8moTMLxQR/lSoj7zaz/Dyxb9PgYj
SMBjlf1ha6D277+m57QTJ3tgzAw9eF/Pt7Lay9VXOwZ6c/j4nuaz5W+/hmgPAt7ha8sPF9ZFQNgE
EBpkO4plnIior+uhIix2lEzsSMHKMezLOTVf1zJbToSsV+IkWRvf47/Ytydnqc5eA1LzmFRyqZy2
6QjExPtYrU379HU5/OrEXBhnRUTXpyH3C/Raq+tuUj+Ei1f/OVDtn0BmmGDWHfVJKJcal4ayGsMp
yzy0inyUvkSPyqI2MY+/co5NYmOhJfX6r7Yo2Cekwf5AF+4Z5wjyVlDpRxA/tXKWuXXGlMd8rMxe
nX8gV4zg6i5bFPehmiFrmEB6vG4FMnigt96A15xHLQgYKm+NcYydkgZw/H/v36cEZAu7mmT9wt0a
FG+N2Toqbqv18jQ1GZv5WdHPnDUuhzUH2j07TrdUXBLkUfxsfcSdE5mDbiryrtaVmLAKmLM4OP8r
6xfNkk2NrhedP7CrRGyt8orVNdrqhF5ReQD+sSjMrlvW5bF8N7Y52RioQ4oCYzCn1sztJyxAhuQX
JMdL6ZmeQNVy4w6n47sp6qw7tpbeIwERlH+Su9cp/snnzXSHAW5/CjMAgfQUeJM/9AG7hFddIFbo
H1guBUazwcn4ijCJqojZvp7iQJ57+aENB7A30vEowCVwUmzdbSbma64Rsw7e4mhDp79nUMBwZwOl
xcpKhqUStsLXrqXrr08KfFpQAmdGMv/MJpf/ruuK+lpp4KfBYHhaAjtU9BhAHD5sTDNsoQegqAFc
08ah204nYqE/NRtqxOYBc4FrWNw3UgHtsvi9kjAxebhWFuH5Owwb6swh1h9LS5aqWLAUWlcCBQ6C
uRv/Ep6lgSZ1JX7P70dUCO9aqQHrkzGPEilprnJ4qKz+DxF4IaHtr4GcS9oCCU/nMnvQOg+sd8Ah
17l2zhVl0lbgCUbU2UGnLk54JT3+7bC16EdriWVEaoIHZsMToNU7nQuTRwDfR4DQD+HGWzgjjQlc
JsfSDal7xk/1T0g5SgXuF/DuJpmXeNenvqjkfPQ7mrc0RfAzWynZ4Otp/mb/05PYQLG3/todT6TZ
cVnGyd78Skr00/QXoIw3r+7wAEuA2BDZghaWM4wbOOKFgmRpsWhu9oULrbF/d6k7zwk93nxghj62
c9+QYVIXb3Qt4ncVrUa6XMIgdPygJ6UUYrYt511CFcAux7KF1Tm6LFifc+gmH74VyxfxuR0wLo3j
2UDp6vEXjiM+QMKBGyxMrUG3cfmTHcyAUULOKh/9RaFQhrABGSvrw+LIhZ6xVNWTLvSBI7uzrHdg
BEstli+upCmWavWY9yPlevz6WrEnkM4Ze4PrwCU6HilXPJBN2/AUQiF5U+J+YaLBJIyeee6Ohqg+
e6iYOkp9iUiMN8Z6Pk2eKpzu66UyIi3YygL8GTahfrVK+qu64+xxlMFg2IEtDpOsFYwLeXiViywL
nRKFW5DZYXYJhU9MQVYuYsNM0FOd/CpaxEFsso/MR1ZzR0j3Td9F+fUVj52zoGWSneomRWg1QVEc
bbEKV/HYel2VVOFKntKVj7h8rrGPCiIBEP2TlRn/wF+w5swVy0Akm65GSz3/EfCiBA1x+g/Kdxt5
nBJJRtEf+8cK1EqTFmiOlUflGGlb2aaUHioYdd7eZLkJTs07WjNZFLmwj+LBZE9rha3iSbUjG9Ix
on9q4BJdPE4lDsHaMR4xRL0Z+hjy6Pj9IkAPsk3h5IA/JhBDGlq3nRaGHh83m18Cmagn/nejLeOP
pa5VSE84ThwD2dC/WFXghFf8dKFaCGocr5XruFAGtMaUVSQse4aOIf6+aKghH8gtwlH00l/h+sDz
H5R6dOeXRtRR1ehoCIyEAvS1lrfZhyC1cqPl1sBtD39DYvd5HSpr2zowr+h/QC2iOslak1vrx4ss
gp2BEeTTBoUiTOGaj0IZSlTSDjnrDSyr33MmyHXuF6MjLsNu43QZ/cqcSCdmQuyr/6yNMEBBgzvZ
7C9D9XJ8XcpLrZR5cVCgV0V9wb+LxBEXTKLH9WJ/qjWy2jzS/R1LRadAGzO64lJQm6UE8QaRy5d7
M89GwP3TnYWu2xfJ3x4NFFkVJVsA0yD+MNMOF7Om2McobA6zsSbWkRrDunDOFmwpPuMZSh65aJt9
zsC/4j6cxB044YvYvfAd7TuK0WmWP6k8iN987OkT3zaEl1IwlfKgwBggjNvNlFX+2CXUNWrIYZYE
RqRPXpgs97LEO3G3K2/mSbF8J/QSZ/RnDLVyQfW5qif+rFN3AFKAsC/cOc4cg5/svrQwckYsOaX4
XKsYb92rsCBievfFWFlLiUQOBYrEBEeEVWWWMIDa4f46JIG4o9Zd0sjVvKTL7kHQj05+njewbtTQ
7FWFhp8MCkeSFeduUR2odLmVR73bGhaxRkI4KAGkrolVewIH7EAqi1H0Cwr708cCNklnoeupxKtA
GhjyUylLa6rqRCYkFe9VAp1bV1H/rSwgUMkgSmUO7moaNSG0MtzbxTkotSeDLvlB3WPLVh/mA87N
eA4JxAK5fDzD5l0by2OVaVMQy3VIJzS8MQj0LDP+aLwSA+wJ7rfGPFrJtEs2RLrqqGJ32ViKFT3l
5NWLnU+ocXdOjc0ge0XNNX0OieVCfJey6I0nzQb4EW400lxj30BusK+SdubB2WeWBBywb1JfX9hs
/WhIlgPWyAbKKtSTFcpjXUm2sD5zpklW08bKAt++pD19VxAzsC5ImlyTB76UYnjdF4dS3XGFtq1+
4KNvxO4ZAk9pK03pWzZKF6umhyNzQo0qMMS9rkpcaBkAVHhF7g1jMolgyQS2NXvUzzpdz2ALNTa+
ZfN+QpkClCCg1jANUfEp/ga1LXip+drxZlWKsMDuxlmoAlFff905qqojJNq85tQ5Qcf3PXUHI0xe
iO3Hv4SMyRFbWDA+ycvlxU22CsusyIzIVUPnWBBQ/g8A+ZShYn5ikKExE1bOSTVQbhBkQ0yERyPC
k3SBusUdsIPntI4Bt0ZpiDNKfSrxJOCwftVuGhSwzljDdQyjVSk2IAbkrTdqgPRVwoDoOgx/r/OL
Sn9LDOv7RfjqUJH6Hj8wEaHJLPIFa4gzSEK8Ls3DVKpd4h6KNWPT0hwVn6pAVHglI2ymU55SSWM3
G4rEjEIvgitnC0zGjtY9InXarXTgcNlnZyzTexnN4JoN53UsFagC4EBJ3d9CyLTfwFlltVnw3uNq
L0F4IBdHlzAlBbEw1zIApfTlWFr+d+GG38CcLMj6FYbTxvxxhtyCJQlYfAYZH0dBUBQHp/VO202I
2NopCShK9NxaNc4KzH134ysmux9a2FX5s1Hh4v6lUgyuhtIMlU9vQDWdNWeYY+MPSPgOCnu8n2Jr
a/R/wRW7ux9eAsz4lRCFwMOn/CjjRiUokjUoTp4k1cUOmpZRcQh9u/RtvO4HL+SJjLPmNHTjZ5MX
DOon6Qt8oCTerJE8ncEBKE7pGoh+2jTM+xrUGNU9TT98b8qbVeF2CwjYcjngLPrz2elwabbhh+Rt
dsvzb7+pT0tqqk0m+cyvXsJSr74TVkl5AwqdwQ9+qiGVdTM1BwuNwd2ZJbMHbRViWUO9hMWdLqr5
l9BKSTuTNjy1vm4jfHIqcX8fPga6EWQiS/O8nyCTkeqhWftMb+79n+dy1OZJs+5LlVX72XaotLVY
PnweOyHyf3rI45TZI4V/rEgJGiEhxhK9HWDRCmXa/IJO8/+y2VoK4HCyZkTweHV1hZxZFWsvyLJ0
6RwO67z/KmC6kqWFg9lp64915BDNhZ8p4duSOE0t4rz/PNYj8KCo2McVCsfjDzrlIg9voKL6l3Z4
QFT/UWH6YQAO0iueh1jEZbNC6G0Ps/TwrAadO1RyODSNNCTU0CsVRsFRmmDYNDHCXEp+Z1W6avnO
ifEZiFOVjqcgMCIr3tc0IMxWb3zoBwEzrvM0YdGr3UY+fQeGcR1hN7XcJM/sgPpQkbuVmyv2zH7j
FAPVHiuqLHgOj1l36VAEnbaR6M8FCUqJEUHiwgokIfa010TFRqH+w+a/kU87Pza0h0XhjfIsrRzw
GCzqCY/BVUzcbvIW2QUTeOYfHcQ8RPdEFbWf4PzMLf9ju4EGmtqXgeTl0ijhjyPE9AkOrvFVm4/C
Lcbfm7VRx3L91IWsOCYc5NYvmP+QCYLP/2IyHEDmnDnHEh1JI9VOUgziLt3h4C31BVgZSCa67gJ6
aRmktybkSyzaOaqKcmvFPlNsnXOMxaOTfFjCXMLb3mbHEfErGlL0KJnoTvTSSAo/p0NOQSFBswV5
fiE+wGx4tFcSvtWcazBDBNU3dN25QsLL1tB1uPrW5J57EC/+6lErYXWUko5+bTYTbX0qR+ulLuMC
TuT8hZ6TRHRnf5pda8xeOAUqnSR0zpsnTTlqssy+wqcPiRYz0jALk/YdL+wBFD0MUxk0tVMeWbI1
3vPvEi1cJmShYe9thndfHzFCNqU2kqx6n25xcblhIa95x1BddUELp+9Dpl9coC9GTZ4QP8/t1j77
3H5XVkwTOBjSsO4IeDzmizKqzB3qfjHoiOiLpJeyQE8GgY38Nc3lYrJadDD0Nk5lsdId3ORTmdph
QmFURgyd+pUNlh7YwCz/MypebJ/ODhjcTeMA2gXZGMnRT2p+Hh7+iLkS33tTAXB3ivOPj4vVZH37
X0ddNJLJHwGg8+cEo7c08llliaLM2lpGxzr0AP6NzcS+Do48k21XJC+A5fUGORnd3gEC0dh7TfAI
gxfl2VuTTXNbty86HL9ZeyHwfpeumUgw4qqWi0W8xfo5Q6NcU1CNVDYRlBpml82HgEch8TszQ1lp
GRPLsx9rLGp2q7NjpLtKPPNjglsY16jzX6faSxvs4/rH/PPF7Ntox0GcNw8AJ2zaSemX8jCBQYJb
JbT58j0ARTdwrC4mxtjR9tBaa3DzHOz5+R42JXwwQPgxrDRkyJg3jp5LmLFiC04DH4AkHOIXz7mv
JeYZZsihVPg4BdPuALth898NYEiKwIGUlnnvG42PQ+Z/YlF5N9idA3CWRB16Pkk0KbhVPIekuaJ/
olg/NeuqJigcQRP65ZA2TTEw5d014jRda1jV+nbIGfpszUPUJLx8TjqYMZhhc9h5Z8bhVUDnXlxc
/hu30cQ3aAKaydC4Nt6pw5af7pCrx8AIhsScWRIvROx8j+stBoT2dYiRWxY4MkS7KFmgPuxUArrI
zVDR7GnRw5+FUaNifz+dbsiyof2bz2cMleh4XFEdzDQh4RtUA2vXh8dzp9sADRHqEXBxN3FM/rWP
g6JjpyFlCRn0XuGzO9YFp/n5N52gHWG7/Yj6E45dDqOi6azmk318GXE9/6sdNi3qKeXv05Jrw3e/
rRhRIlMCNsQFwQRt7/kf3/bI1qwFsnRsH98DJ6H5KaXt18rMkFC/bptaXFKOK96y1UxHkBi4l5rf
nFxK67B8chr9GOlwHKA2O1I+3+cG3MxFVSHHksympQSCvKf1cRhXGkjs4adnraRHA9uQho5CkK2P
x+4Rc+g5Ux1IcqfPRszNYWWKWtLHt33InsuxdOY110O2zyVe0CfqsybQW/9wHkeDfgablbBLb7TW
ZiihZji+d1MjOkvcNDKVjmwOeBpZLwkiL7gHMej9s2LDRGd92HaWm2LI5EslJ4581w1LNKQ/vIpV
W33iXZ6OBs9YGyRjzcE5zQOIGyf3TU1N7NjCq0hql/ehA3J+3YPl96DhpKDuzr4y8fl3FjZDIhO3
D/55cUJrRTO5SujBTVbyTzUiD3aqDO+CTpP2uj5RxAQtteaMpnwUVes0w5Fv19p+air3l1a4kO+3
3bEPnDpusQa7UQJ4yeemvMk0IqdMFdECpmoA1bV6QS3KOtoLYphljsZKTdSSX5QCyH4OVLJeLtMO
YJjaKvvkKq75PRie5/rfcevC0tgDraEgUtjmPkw/Q8BJqoAmcjehNE6UyGhg7ARxXQA0j+G1o6tt
CBzkta5UG3QS31XCdKwrwREa1XDPRJMNo7LCGPEC3kjBLTyDKqLcaRcuqSk32NX1cvQihXG0ocaX
0fQN5JonPFuBMT3MHiASpNQS2sLsq99QazU5TRbNYoGz7jK1IOuvfUFFF5YfJDKkG0Rul9RQf0j3
AqocccTZBENd2z6xcdttyCY5CD/1aJOtx5GQp0VvR4PC094IEnRFc8ljqQiflvRjqrX9ORS2W5KK
jsTjmvVJreA5BYBFDpOWji30cp0d5XqSy8FDZU2r9l/zfjR8NGDBeqlq1LryW39zvU18fREao5jt
Oq1T9x0pWfD/mPNzbKaonJZ06WybbQ5w6zpU1GVEmljbcsU9YvDFQB6x1wGCfCvi9EsN5rWpJ8VK
2vbX2L2wsuK8l/5fcrdaTg2uWx/+GNgtyB9WHgoc+87sK0u7HfdmwrKdNyVS/ddfYEMYpw5gYeOy
eenATlSdmOKMwKpG7Chz0jSAH7ad/COod75pA3iHmKGQ/R8iVmAiJpO54zXs4IlIycEDIHu8pYor
AVj4q9wW1Qxd046KmctysDQr3Bqv/7TwtcbvlqOxWDxV3vcaMMzMYKN0FYL/a9pqsJ/lzEKf9d7K
4DnTyagAPZc7Y+85HNQ/KH15pWT00ggtwADGPqx4miZNiDzxefuL9LVZX/ChVoPVLF5dNFHh4LQT
ryF/6mtszKP9jLAXF+qL17AW4IChVWw4EkspNPOO/JduLLA3ycQ5wNv/uiZhyXRJNJ6NZlehDcbJ
/MxTObH7LCQ8p5QCkMElzi9dK8MzM0EBMZPa5EeoHG6zytsATcU9RkkxwFwzjHWThonU8WvSWhD8
aSv8ttl5l2VHMWSsYb/f8xBQG1EI0U0uny4O0d/vnimcAh5Si9SSC3lGZNcWYWkG0CXBrkLWroZ0
T1dRs9M8u/R1X4Dbm6dDTipQrpfp3ZiU5mJZQA95/0t9Roo8qxs5KDvoZTNDwMgwkIdMTTj6oX4l
BWHpj7lP6rGvk2mW9FPl9eX2d9KfK5N3jLNZJHPm9YQdZp42dXt3EQPOZ9lOQBiY9jDBP1h3g5OV
UHtWecCQY4rJEDZmGCrnyacSjUOKyUdhHj95S9pHAVb4zLQIuVGBnmJr+h9Lmf0ixpXm7zZSkb+u
ocxJUBx9jiNjJPDCyPpRSzxCmXtuD6Agv8MKWFSfNwbKrAne2lPp8OCqj3f+Mbsir+6XsQecNA7u
bpyfgD6sn+k5GJamAJ9EtFAn2M6d91mWcqjDZzqSqm8hqL+7vO9L5ZfVJ4K2UWLJM+d+VKGEXurC
lYpl9CXabvYQlQSgNZ9mDC/mDPJMUutQqDL0NqckTAypg8twD2wb/9Jhp/zVfNTo1TOH+XUHGDkT
eb2DEWmfy2b3QTGiIKAaLylaaVzKEEUcVB1PhUwMQj/2Vb3TBC0B1KcAJe9wl8jHHUiALfpdQE+4
iYoX5Y/oulR7hT8VxcuNjF6XZQbuCOtXe9DPcvzuv03PNHf9pkowqYnKqDRxylgdxR8SDkROwh+v
ziAZ9nvIlgf5VrM3PKMcUlkjYcNLAXAmld+4i4jt32U1bYSYQr9C3y+w7ZyDVyoHfmBdtXyXTrbC
CiUjfU375cCdU6hDXoXndwfItuMc6RDRbUUuR7wbLxxhSab1Y3RIRUYOMnrPSHw6Yo+K1rVf7N6C
M36m3HFG8qBjfDsK7SeK9xL86bpXlnMrXQ49bLrGmjMEQUdnB4mpq8MfwLzGNDVUf06apuJxX0OU
F8XGSkcD10yL5y1UiFAdwgulNkRwM5yJLZk6KJ30qh1ilXZhwCVZI1SYPl7JlWJoRuD8LYSTFL3e
Uq1mosmwOiV5n3LPT5UU3n20+lHVfqm8HMPi8y3IPc1opOFd06B4b/AM0jrw5mPp/VzeCL+GHcGV
PMv+ifUGzz3jJuM4QhsxdYzNRN61fgim2MPQEJZwiFgrYBd914ekcifqxXlHo5oeaZk742kDN4ys
rWdpla2qAOOA1khfKpWhb//PCB9nol+/DepyQMM9nynECBx6oKCAklepVUHZrdjjbZTEVuhdnWO+
NfdAo+WZ2HfOln5sEGP66O259OTx5uPS1MrUnfYnmsBwrfrc1ZCaIliIIpBgwyUooTLnTim/BDTE
XEFu790IKO8CunF6X+RHQqK4hkVeelh2YKOx0yQu+92f9fPKgY0vTvT7qp5ciKzhplcWFIXevlnt
u9OjtlqIJYn36s53uCzmV4t7t8Ssaky1YQ5rjUXFk7YE7sAUfBxtx4krXdUiylI3CFCD4WJACdvH
ahm0ixN0Fc/VOpd/ffeQEHgYdceVFrfbXJZGgeL+hCgjaztSDXHO+u6YsvTL2CW8XOjxry+CHeL/
igGkRitnATEohDaq75vAKVzSf+p8cQKFZwnUPxIMZuVT6CY1F3kVKJGtCMOOSkinZ7NAZ5sDQNuK
SiZlM2R9lCQD5Z+e/p9GwG46tS/9J2YQ2zWluZs6jGqQ6n4nY4NHysDIMcta0ih7UdI2WnXHr189
ohVmMjNOCgXr7ghFZUt2+zS0XlQmieRBRJSvvuIkhlJq5jCcshk4x74StecC4gJTbJlL4y5Kbufw
mAE4//ZatBAp7tj2OY6rE4qXMXrSZn/4kWZVFUvpuOfbKWeQtZRfhnvSXvjHa85zfT+omA9Ggn0w
FDOKgxYx6rfGpPfuaxIa5yUXugZKGog9ai/7AD9OBF8BIOFeXXKlWM3JKR+Dt48+PV8Te5S7ir/u
9L4bhanfHYUdV1q2Tync1I0MV8qEGgylxNu9oZFPzEAazw00NdmGj77T0SpCnm2rkcgQ6ybC9LnN
wgruqDccJgcK3jH5HMfba5mB43/ZCCqVl9qFt3rATnWplHwCtsVSZ4VfC4scbVYQGYdq9svk59wg
RCFe/BDMIun8eJmeFC236R2CATL1l9CsxZ+1nuu+2LANNK90iWebH2dvTG5l+3PwLB2Sf1JT1iyt
9yEE4BcZQxRYA/Abttc6JxZxYpAvUe9+FUPKWF6zzaDwbMsyNO8jIHQLYmDUIrbl3KydiPk4gMXo
I05AHQcZfAJgfNIJLY5AmbUx+R7dMSvIs8OPo4zhC2u3ilSUFn8xdmgm0orKI1osYo8FRiUrvv3k
BOLYhV+caSyabWotdUW9MBsXnQoJu/eNLPUJqhfsKwA5MCzGk+nR9Qy5w1uPJ5uvAIaGWuXkXmGy
oatyPy6ItO6RZycXHn4e9vLRn4L2kUVU797AdAhvPDYqdl9kVC06CazbdfbRloyg8FO6gLzgJQVv
YF9MyVrD6frfnRp9ZdtiIu1TZWBzDzdZwILCOCg9Q04DXDJyD3R65gZb7Kw98r1dHUg10tMnm3Dq
wJ9wJkymCygHGCuuYiE/+329cFAItbhPwqP93yLjyyXwQgZWZeqFKlMRcsnkPuwF7CwCA1ijmLmm
tji5rXjS0fa6kC3O7P+RYzhk5HadrihtJWu0xYqqbGbq/6VCb5/qsImRlSbeWXV08BMFv1Lk3629
+ee7GAH3AEjXS4xZQg1sICnHh6sG/d6LFUZl9VGmUDXZxruHe/FEafmWzBRKEEHg6EuRks9mSF0q
hO6tLnlM2MGLZ9n/4xFge0rBA4LqqOO7mBCXW+63SL7o0Qevx9v2/KHyW4m2O3r06ZmMuHsppHYO
gExwDC1G0usUk3FhgxdmbWZSPnxcm9FfhJiWPbKCYH7oGs/Wl0Ldv4ETvoV1pbiJn2IuTtYrl31I
qIM1TjoxnRP8MIVWEKSH/wt6ZfOxGDn/+9OrCZ6nao+Zj/NW4Qr740gvhhFiWNOCmsFi/Sg9HMS4
pSzAFyRzbGpIm2iY66pCPEq9bOW3IDCJlHEYANFEyRYV28cJpZrFoaSoT6p2IpqmO3I5lsR7y/s3
JvkKiloUCWetIQVRLOkpBP8DLXkY246edsu6OL8K+3wv8ujpmDCZKq4mVkFgD2983E8nOayNDlPB
dGlNK77TwIEkT3dfkx8a1u7ubM3qnRn4WdtuAu5BItCQARYi63kv5ncEJQRMC+wh6CQ2XnW8MAn5
sKAYtPbJwB848ttC5HSzrSD4ys+h9FbqIGg3T6lck85xj1umSnWP5ZJQQJYawK5kFjeosFuOQjyJ
D6khr2pSQMRxSAqZSqFQRChhrzLjPEEaX6ksDy7ZAoPLg9Ld2M+MbKHOHNcB6pVmAz1IkHVoDSo8
dBgVLjBOEAzXTYCc97rjVX6qpIdHF33aKp6kqEZ7Y7UZnGqGvf6BZd1V0XFtzPh4ZWPB9gVYUgbC
437DE3jjk70bBGePqhfMKHkPQwLhruHB3A+lB+YiAEUA7P+IEti886h4aXYGRh2Jp/RUEUxihrTN
RPTrPyg8Wn6zl5M6r0SBeiPTj4xEuaTaHxWA5T6YWyRsBoV8uGUrQWhZdEyd+7wl3TFDOy6pGcJ1
3lG4LG8ryxYOH/JiQhsv5+/R287Yfh3LeLM/K59bYtf9UEhRxatcV+PzK8HUS8I2a0urkrIKC5sj
4GIatDNIvnF33ioFV7c1kjKkYB2PLDFRy+OaCSn5jUXh4oxGVZNaY/MOvHw0/aJ0GnmM5r21n5rz
P74yJnp3uTi1BtTau78SyyM5Yhc5ujqkUPuT4eOqbnXrsh2XyWSmtIW9TSFprYJcUMq2+DHjcE07
XEdu+X28jOlx4EuLK3827+8L/ARnmeySi9/mFdW36tf/ksCNiWY4AAtECHrgO1AWFuONI2a/v6/b
oJtakkjeTHh9v4Vq5b0pCRJgOmYJXh85+zDzGfg1ECcFqtuaxQsQaT6GLT1yxFOhpvj60OEZro/7
KSK6vh/AoVmmXeog4MhLSt6amrByREC5dfPWqoqXaqoffGMnEwWb+2sxOCrFiIt77ZWWi67HfO0y
InUGy2lC0a2eKVgXjZ8p/DsotCNFilx8wKEtFf/vA9o+MWCbQOLRcggx3dLv/dbTD79rP1GsSMx6
XzJQRONE4vEWadHugH3TzhKYm4m8NVZneupYA7LwEq/hcAMLLcvZwcxELl5XMIkl8BQ/4xzCrSyl
CbHN/Mxd18tA/7bTtYuSU0Gkry+MoLUt9+XYUJOLJHW8g4sbcXBhWbA4yNa0QJi2FKbpALq4Ti+X
McfqMpznyd2QOHeVfWYuc4ADlt36yEJoRGcfyieKLCTnCvjPXTZrqZo+q0/CXtVoCqNwPPutmf0E
35dBv2DzP19ae5X28g8SaOKAwudd2zmI1/XSXwPPACaxcINhPlpDByv6OAo1AvixEGWBGS2RNw+y
v1wTcVPalSt5pBSLqKs2t/6WzQVxO4bs5SYDsl2mu/od0tcQ2BpjHB928O8RwqFJ6lSR3hR/rpuQ
YM+HBmOwz5ja7cP+RFm4PEbKnQM96GYyA3brcCa5Y59+wkIT1blsEir1ByzfJ7dn3/2a8FvE+nCS
z7aSEkGYl8EWoLL4Yqfmr/9m/zDhgKuxYVnzMr6gKKahfIEXtKRE5Rkg+SaPVMDAu6AYJORabnXI
JnAyRvrEVaTo/+NHVYBb1vT1LP/4tpF/F5cGfr6c+DEoRJkYsQN81WK4X1DehHKurgaJLJERZe//
rZHmdh3ghti0luRwXm6kdBUINWJQqFl/YfZUrI+amLPv/1ulOmPchR6hHcnTGZehCioox2wAsLR1
dm6LZb4ZNN3JRpwz82ZDioGwsVXf1u3UWV/gjGULd4o70XT73v6Fkxm2Wbc4CCfV0PBzVBa7gxPm
7xwhSEGtOpn+RGvZz0CdCFu04bAKEzAzSQo/HXZcAM0KQ6++LhEnRM6OfMIa40mqDXw+6548UYlG
r7BQfxFoo//2v48HQxFqAHzTQ8cJkACy1Qf1cIjfPsrCROf+DZv0FuIsMWA7PJKy3ZmK22elEmyE
y6wFmQTQFJikJmYCFQs8sLYXTYwpkfkzHGLBOvI/q4Nyc69zvyLCASslGU8VH5z3vegGjOHR9fUZ
016v/hrDpUY1UzRlJitCK4X0IsYutgw9vnKzmvQoo0vvppHaE9Mg9SgNSNFsp+19y/MbsrMr/rIF
MBRoyjc5lL9DCzdBnALdDXOQgV5nGSXLcgW9DgcvG2tt+tNT+K1IGmFDmWQgmztG9fAAcLgSxIpa
Fr9a/E1W3y7kP+axc7ckExHNBo+vuhqK6AduXJnNVQ9H9NBX6QU0ZXE2IPus5rPzQoDcRJDB+6SH
L9bXwy+ZJ8VGmvodiXy2Vv3K2+HFlaYjwUk1hB7NQM1Q9fUGW0CChTy9Zn1EluyGXlMR6EEZrmSc
vmAVqVtx1sJD3R5hRCxfBUgA7lfKTnnTvYQFlcwHdu81HMEXhAL355T9kWWij4TP5dL/+OA55t84
mfw3bfuCwh4qgrV8xjuHQd9FRhKiHGYW+mvzVBI36pFNC/L9F1EBWh2BNkyR08V2yqh4NPTNB21v
eyI7k9Y8siWaEd2/w9NM6v48qAwVx+vhXSkc0L1VzdWesOc+1MugQFpV3fVIYok70hYfC63iWQAz
l/bcGUE5LZPhFVxI/jIMekHQrFJ5vYyGxP/60EIcd/5HvxXvGuoVVdEv+8ZgpbeqhsbhWJXMDjgW
CSK4dDrgwbcb9yF4DJHmRAgA7nBhv9m8bFYeQdWZcIX0HdP0VR0I2o6/ZuPP+aGwWH33zYq5e53x
NKg9XLNfQeMeW073THyzDCXlVBr/SwJ8pQhT+WHsTbOTADPsBfBll5Leo4nOFaIZn/E9IBLsRJP7
b1wABo2W10SnqYW0bBIc+tJLYc3C1K7vATQkjwCwUrcMwlg8j3XoW/FQpZuv6ILBm06rpAnAKuz5
qDDwynPfxy8xSzSYNmmNj/ZdyQxogSnbgViPyCwaCa3BQgtBGOp3gXVKU+TnvOvsgYarGFfZeMEr
G8a7d11m1TUfOCmS6sXpB9kJiu/Si9ZZ4hVH7iJVtHHS0j4Yp6fMmO01eYMoDb1qKtWXcc8dDwUX
JHENoq5eAkmA8tJuNOZBvicXY66KJSj7ThoqQRIXVX7oUYEKHBpqeqly7X9Aa/nB5QIPAbY9Hmub
R+FMZUCHW98d2lrgbJUAVMDGhDaHbZHeQ1BiJXQG+x8GHgJFtIjwQR5Lpzr4BOqvEBhtUVigbAAj
uhHbxK/9NxkZjmVqK/Wc5NJk9pt8o6Mn6RT2CNTJFs21othtlYV4sEj9eu5RCcTjTRkEAPqCQ4Qi
pqDUd/vmIh/9e+B6tgdRY8V4WB7Mz7GHswR18sPq+po75bYpXm8FFzwY6ts5xaE+gtI+NGW3PTHZ
30zBwHrpgE+nGSiIkmY5AUVl/Myw5Bc11fEr777mK+/esC9+SlqyYfMEbZEjg3wKWjV9aFDB1P2C
PbSYQn7SJzBDj7Cd4asAD2UYBr5A9cjN/PMZ49vAfEyQf1ryeeyK4xb7+e6a6oFq4QPp0ygfQXti
SDoLMZ3FdDWVbsZxfZeGFL3H+rdmp+5oNPkQg0Rd4u0ut2fSmyAVEj///sy2ZytaILbWXs0fB8AS
Ew1Atv2tSwpMEewUMJrLFSsrSREqJ3pxsJyONoThF11pBXunm4fBXLBELaVUy2UrWcAzs2JTKJTL
OJajhwQ1/mW3eZvWZNCye20X9lLCXRaD4flEzI94eFh74qSPXvqfkUZcFas7talz49hamK3I5eVa
FOutZZJ3lywWuf1GAFv4l7m1DQCpOpyAjoTbzmhs+L8pNe4WlxYCGhkvbHiwwkNskHDlcPu8eMtU
I46iiWI6dPxZFei9/32qSam86VZFEg9nJr65xAyu5MpO9TuAfVXc/R7SQvWxT+cl+/R8IDkoGUNm
M/A1qFH7vd80Voi1ccOpzOLI+Gh+1OGWiliCXGDuRAWXC751sKn25MWwNvBBCBkRFqtcwY0V7YAg
oCNpn9uxLPWV19yBCiwSW0Vzb036/3nZ4YZ1cpGKt6Rkqs+u6AViiJCTXSekiZ6a1HivuDolHP0Q
es8m4GO0ou5fQhltY2+cIFICJ8j1n+FgAePDA/XGV01uD5i1GZuXDTgmxG4PHhLqKXxS89ZmHB+0
DittV/ohWSXIZAK4ZHWvHHFxXv5iO/sZfHWMR+GxXZ/4+tERUy2okYM0FRS07ENEqbpAjWRtYumY
QAkm6Pqqnz5iJC48m5HC9wWEJ8OhosnLq1hpP4AdupGXglcGj49PR93PjouRR1HLx1R9QvD5hMrF
wd0fAbzoQNDA8P0h6thc+GEl4K8RfzrS1nKMG5EDuWsWmd6b4Ju4BsXGNVYr7wzyYocuImEc/l+B
cZ9FvBUsFG+jCBddEo1URcv1ghy6fttjti3hU36UQ1tFViLwUe26Wj3ZzFRJN+8oNPwtDXKZr8fu
IC5TXYeEFYPfgA6wCP25TekYRPTHhkTC+1K0nI4cVioDiwrUXfycDV93+Ie4hdFt8A/DMcnhc5ey
odmxIYORJyOvbFwGDXGefhfGxhF1mtwoFCbkrywHxPPg5t+d50fiaE3FQzMEoh803xPLgm+3hLVz
f9QdPzMf+CQvHjHesIzL86XIpQSz3PhGAO0pyCbVrN5nH/PQMHfTiQ+jhU3N4/Cs6SPiJGDE13oh
TmcbysTObAZnIGJlCRgSjpbcwXv3TNRSM5TtjsjlFXXF8iMcTpKLR9k1/+PASoAiYWMprtqMZRah
Or6pzEyuacqcHmtwEy+YylFz1b4qwGhJ07FuFT2WeL9kIdpbOm8fU/mN24176sAJffpis4sP69JA
qN29Uv1Db0uX2grVdSTPEfT1JuTwjoIE0ium6XXSTBDE5sXMAAOBCPWPuf99bCfPj2sfdSlw/gSo
8QFZKI3D3/0VYHRenZcDepCfJAkgBBdok3l4uT/Y4R6BkTxBA8YJi4ZplhYJzWz7SK8WR7NAej44
hURX1hacLv0K2nVDZqSlurLOHebUjlH2/l08NhTnt64qWHuKddVL+/NjGcMHfQ6qWye/ej7jU2Zz
h/bjRORKnMTl/x6BckZ3XunFLWuhugsr2X1jsv8vaTnWqmzsMdjvWZCgnn6A7yGxpjpTYdCjB4HF
AAdalnFBADilxggcXjDYbwx7a0BRxgubPZ7YpX4ihpuaMIMfNmbf2JFKFDy+Ss1ntACMYnHeOOA2
ln6l+HEsQ6RhJEgXNzlhxNYYObOYWAmvSY4tXowF1xrENP9ox7OP83pgGOQXKtvHE2iq7epluFTK
sDEeKSNJ67OLqTzoqRFUu0tY/7WYNn/4QKpfyVo75zUEh4I7eHJjuqtK+m1AMVQeVwxbHd8R8t2j
FSvzmoKg1/NeqhQtHmGQ8H6RAAW81MpINiwvC6q0wKJMM3zoTB3xgLitqik1P17Z9jUHLespHYza
tdTHSgsuaILNbnt1ugfF/I+egvhPXApMKwRiczMZTDIx2JH6Cs+91OKcgwnZjFSwFcQAzmYByZZ7
kF382H4DoQyZP4Y2LI4DaqemDLjGKqHy97VnsG6CLh0iAnCqi09XflIbuarxwGOuJ4PGW+i0hHdo
y79y6i2ihPHUUWqFkG3BsdURf1V0RfQIAmf71a9s+ofUVYcoRlPkxq91GxylDZERSYeJajQd2qMy
HjSWRQa9WIYhsBYMDCdCHiLu+ZpUD/28rprspZMI+malA1MvwtUSOncdGeeu7y+NlEougIt+QVhb
NDMGjjONXrc1qmfU+XAOvZnunn8DPFP/UYe2+G3GzTI5Ee7zSrVwbPouyhSmiggjOANmZHy3HDO0
Xx6YnHWen2D1IZ53UZaU4N5USrKs10Aw+zHZBmXKVwVgZM4EUzb4UTdye/N4yEIVDDZL+rBlMTnB
G+WKc1h/AUy/p/RQ07Ttgo55hyzWCn8wXXThlzKumju0umNZMqvzsG0K+FWlv0wSQhGAtXuF/YMc
ADBk/+8mnflDqzkztPkSozc/ibGNkdi5CbSEptfZfehFya1nX2/Aa/26xMDklgcg9DTdnRPssKT4
+8EUcttXwogRLDzQAC5ULiiBZ+CG9/RRcTWkE7Pt8Us9IdXRBN9s3TunlOV7ot0C4da8BdzADnl2
/svZWnbri1bzVUTaobH5ycNarnM55aWGTADwhvkp+17dFMwLQzUz42D2kd2KcfI9pdq5VBaskuQA
2HGcfuW+GvSbhbFztt6LcnRdZPbMFLQOk9Jnn7pSvJ09KAVH0juHp1nG3A0khPqFF9Ar7iathIjD
Wz/I1UG5CTfbvzl7+TCEZj1fgOzMYhI3oJnaLGWOFYrL4jGq9o1S2aqdREajr2lWmsUelC68FjTs
4GMKRR2qGKSnDA27WGCgpzYtzvyaOrGRhrDcei5Kv/65A5qFdwCGud9vYDtDtHelnowVmn14RLdB
8ufLbRKezLZiDAUZ4HevTGpI6tnP5dRxtNFYl25TFjljj1c/qsU5SWQ1K+Vtedqga+Mccn/fTkfs
UwBcaTIx/A1IjCxbUe8ZTEm5G+ZnFz3fnJcTWw7hxkr7cZ7tsgtXsGYkWOmZQdLqZ4VcN1aHtP2c
8wbRpuLqQzHpPF7e2yXAk4tJ+fUBoebhhRT6R5hi0BGNPaejLm58ESDb0bQTU1nI0j3An/aYlk2w
uV60KLivTmtlt8Y63SEqv1mA9sU3AXZAVdiZqdda+qo6Fu9/R5Boom3M95UdJEKYacOm3IzqNm4U
cYglhUFPQk06QF0+Sdz5AYJEuJNAjHhKDpSG536vVZkS/VTPty+BVeG5iMUSQZGFuarGJ/9PD9vm
//C4uUiaNOgnI2roLxyJON96rBKk6+Pv68eWQYVhaYBhE6ZjVhhffJc6dFS7r+K5IwWOYz4CJgFP
5RGgWpTXNyA6Emp6piflBW3t/tomIWd2RFTXUYoBlXRzlHgS+WXxqXaEyPd8hphrYbA3CcmgkjPu
5l3L6+UoJ6vHehEw9Xp0FFW1Jq6LKUaFzoGmS+0PSgo08NxT9VftCrFSOksgAONuyvepyS6Bq3Eb
8seFgafpq3Nio+SnzloBZHKWApPlRBVZhRlGLapxaZmhy0yBlej7TLqZz+BIzH4/4/CcB+2IKID9
Yple/W5IKSjQkhD3vx4lvXmEbH4V3EFZku3Wga6AbiqFcln0Kk/FfgftBDK3J40MZmyJwK9FPHdh
93ikJLbiRgGRb+QyAeJpOpDBPySiVn2RxWYuN3ECv9SpQmdhnvv9QDkE/nRik+Q2R/jzbMeN4mwX
Ss01qetXphF7u0QSKUf6k1XsYTRFqTFXxpQI+C4Narq+pG/KNli6vkJmXCMwO99lWbUNuwNhNgDm
V8CvudkY4wQAqFGuhVQZFQiY450pmpGQlUyOzdwD8yXp3exqazcd9LIMkxdQjFH0U6IgzZQ1lBGy
Zot2DzwNKbr/3nlWOVx6GkaPLcE+h/1TRC4rWleM98q3vZJUZm7YyEEqYJR/LJf+Em3AApN3lSGG
ygyFvrzwP4KI+X7GHpDc4hq22U+2mG4WwT1B3btLz1YF6FZ+uZE6DK3trKjZMCPUiGcwleNaRNb4
mJRP6scylejx+wyin6jq2dgDOg+OvlBX97ooBOcOh24Z+Ave0eBc31YtjYPMG8dkfyCGz880Sqt/
p4P/pKDx+V/l7dP2f7NhXc2fMs6aKfioA2PqEIafHiuMo9cWma+Cx3KPU4JGUC/CbeIiKBFmrqk1
F9y48X8hZL6gNDG5gF6OknYlkAq+xNICoa72+5tqz4AMOoctF43CKzFrftNG3oeJcG0eN8VYUo8C
d0I2kwLgU6hkZQBdZS/VQs/ncAvwq67GIj84TPjfT86Ywpbzj9sqNF1daoT9Vd3aZd0c04ozeAVC
GaB17K2WIHZE/i9lzkE/9n22Pfk1chIE5+CgBHDpLo15OCJOPT38nUP2enCmTZVONYyIQTDHctHZ
rmnc7tv8q6MDH1+04opbVsGASQN1/9Fa5wPgCEyaqmK5XQ1dhBcKJHafRh2s6ZnjvGh0zgz8bOSY
zf5a3nKDHacXCHazDtMRi++MN4HGnwiCQZM/pn+Vfct0YgFMfI4Hn9kkIzcqoi22k9heUb0lHs8F
F6XyfA4V/pKvsrBHjclGrQNy8/Xj4VUA7RLnW8/H6AaKknPXgYpisQOQsnHstn5uGXnbdnKcFCmE
HsrG1hl0yeB6LaS1g5bGQIeinR2NcN63mfT/W39TopewydxL/4YFFwM25l/b6vny6QogcvEBq9qh
/h9itwFoit/kleN7yYkBD05RozvXi+acludWkVT8tRf7zmoJb9lPofTc77RqfUS8m2LJxMkc5T06
T1bG5sQL7pNTNwb0AiqpktKQVEupFQaUNlFxXpwsNF+J7CTc38eTQ3gt8ucwS8SmrrXEl6x8qjb5
iW+mArgwOJuwoa4KpviOJqNqCkAxBVTsldXWEcyDx5VKf/kupuhtZxgA39MnoBwIZIw72SRf1eia
WBl7apEHxv45aHpclZ1UwdEQykl6NrGUWAlh5uZpnOBz1vYrXY05wQGa9IHkj8CRhGSRZ48JC/HD
ZI1prQXXI15W/VxBwoG0ERoAmcLFBXc1bEWCvYxy8NVPLJS8DdadtlfhxBr42gH4XGrblKmG9wJ3
w82p4M8tXnzDAL72rLo2AdRAcn+7Cld4UnzuCrJxrEnWC+iFbvYBEVGPijUt51nrJHFf2FNsKI0G
AAv3k/CfqDBlNayT75nlbbnHz+PleubUnMKKY2VuQLJ1H/rqvctqgPF1pzkAB4L9kCf/JE9aczSl
g+nGkiyM6Qz02DlovOVo+bzot1PVfVk3It+KQ1hKFiJQxPEMS+CBVliHqoAxtSoMyacvq/p4M4e5
yOaEqlZOqVZX70puBZxvas5x2eCmwEW4iqVw6Tregba/vIvwXOGeOuCFkbintuGbCzVVuXFz5fHQ
6zyECaG0J8ljdqfh34kNawHJPsRPjLWTjEbuoIpPhjRF6nbBTAz12CUlmRceA1Blbx/tq4ix7ZoK
ghnJLB7i0NWSnzTxIDgeQO5SV24/Hy4eQkM+mU2t4twAXBtHoRzVxGBi507D71X9vzzezPo7m/xc
l8U367USfFm6+nYuuGVIvtGv4Bvw0yJYIGPOdSHNvzVU6dLAvXoQBqf7C1xEmFCA7/DqlmcR7wR0
EFjP1j5h5AwNj6VxCG+gliPX7SQQYGi5gdVYd9bg+hWD94KWHFQ63smVBjAWvozS8qCxFB/V9wXf
NQhNfaSUzrj8Dx5UWJq2mX2ojudup4bxccvOWNQKGpH1hEq7briHNo3+sz/mSsuDMR+R3xx+KZl+
K9H01WrmUyOTM4C5G8eLsEuntqabH7ySo2qarrSktxfD2wvMZ7+n6AWlBBmAcKM/IQ/NPDmYy8lQ
QD//DC9+jDoxxgEn1kLnjKMEZC0SkDyHYAz1MqzowBhZp2VA1RM4Ji8Bb6jEgGE0k4KtPKlJ+5qX
ePc9NANAjndhEbLB6wSQBORNFRr5LfZoQSnn1pYKiQh4TG2bRKzoo+jqR1ZG8XT8vx9zY7oUOVRa
Xxki4x2S+D1UEhWUFAs3X4DtbEdDOHLLh1OQxt2H6HH09w29TzgJ0Ez5l9swFXqTjC5QthPb2IyH
xr3PEKnljt/l3JN3aXUgVj0s/B6GnZ4ettB2SAK2bLO5L2dsHEN1fZb8XGL9ZF7rbcWCBOO3iegt
am+JnkljHg3DNWrI9Yg5QH+2uksUZb2kD2aCxIHfdN9S4gO+4Y/+EPRnr82pAyGp/tLjJd8YNyOE
agvZdYg+gFx3WaKmQnRPQs9lbLMzJYa1LVYb1PX7GYCKRbkUnmo6vY8vDrCrN31Ox5XkCz7xTcYG
NvUi17HcLj/LagDTtEUaWFl/Zx13OZWpiK+808yFXoNCmElZ35FvSDntxhCrgMr4qQINiayYWt53
oooJfnMUtazo1Tt11ixEhxBuSG3jNevzNByrN1ZESucphv/bSghpOhPQg+O9yEomzqIwaflyGIaE
ZMJCl2Z/+ddG5Ennikjum9Gvs6EfWIL3jtky67Y6k8WtR+QSbHk+TRkcXMaqUFhPN+QovqVSHb80
8dpU8UeOx7K5eLEKM1vPWCuaHXqCKNpCtHO1CnjnXl2AaGyMw/yJzgzAXR2ZRQ2DMAaa0VKKLDlq
mM9+FXufNpcHwRmgMq75Qhk3KxYLtUnT9bBwf68B6t57QOP5/Uzm/H3YpQyCpPTIrtfoL07hjemU
BGiUoo9CfO74prRxFSocGwHRGtj7/SL7LWJ0cFzRMfyjymi2tbA/4KPb3tAGtCK4ljReZVUL4p+n
3x91c3vuH8z0u8vMTI2CBRCN4Zd+V8AB/gBcr1ut3Q69sMkD1+4Y3mphAIoq/IUnKN85n6qAQFA4
Qw7qpMP3Mp9IRdv/wl1n+oPUN+OqJEMV/ogzzFVnuQHMqzlljWPkcYC/kQw9rUvx0j4YCZoOJUjB
b0v+Gj3PnDZFqqztAoY53LCuDWakEHrFV2Y1SPfZaBjc3+oDcQhnbHZdmK6vJHpR6ptqxeoXoXkA
GWfgjJyk+fjBs9ukCPYHUmTlS2fWySh0uuVRJFFLfsG6/MKw/c0eHf0VhiAa8bK4cG2uabuXKv57
XCDO01cfili84nuxi3+XnkF5GblsNnGO7/2fvIlkRqYynbETlQazaFv4UyRrTPztjOy8kQzH0VPQ
DALb97C4KpjOGtYf9bwGW1tPZUgRDTtWsp2AVHJpYI+IWQrf5yjF/4b95ruO2uXraCIoyVm6J1Cy
MJO/K5jUgzV80JFh4JYrB6fFPKurWdbi7tIQ/f2kXnLRzwO3sDA5dHRDebnNHYLzz8FqDUzQwTLO
eb9h/SUbHUIh7ZvwNbeKpz/uZy3rzirhPOveTuu2bJrEkXhV0q3PoU04cbPlSuZEEcL1Si5c/a3r
CH10HIKPKsmGWl0uJU/lldw3OoWnhuHq1UqFelUp/7uvUP9f2eT1TY5YGuEWSFClHtM5lhDPxh6W
X8kUdr8UP0F8D0BlJOG+RzddOlWjl+vGPmW8vxugOdDXiFwbdGWfJmnSkpntNeNFezbyG4D2bJ69
Tn9P6zeV7L6uEAM2DBKKvNmZRQ8xwRzWMuUbYegb9ZZaO7Hr4N6nffuipOHPrrHiepQVU2c33xol
UJOwGOAq1WcuQV1mILuQm+PwL4PeUhpGxSjzdJ0opjfFQ4klRuNTgL44BmDqnj8ODAi8dcRdB4mV
mYgrnBsm4fV17vfAW4NEhI3exHIGbc1bLUCA5iC+7I01TdwYWuSmNMCr0UPbr9CiK1pnq+boYIzn
b1Pslgb4KdxQUzKNp79ScE18Pku8vR58+XdxsxsvTitq1oCA6TpJHMRbTe/ssHsGnzTV0eWVrQVH
MezPN6VeLojF2ZUEptPAw7ITPerCQgbsdbJPtPgSvAwo2gsA6XJN99c59ThfPUNz2o3mbnHN+/6g
0Bqm+s4n6I018jUgPw54/tFcOqeXA4Wnts1i55kXc39lpFtZ6n9uYaetiz2eurb+HROAiw87z+Rf
wTjfXRzhGgezzqNZAgMwSV8xMZWmFhBn95hPZMskjyXJ5cZ8LqSEXpqFP78FqydvRpaxMC6PqAm1
BtVqyrw4jQ0Y2nzgAVtLhR9zIfDDj7gviu3nihpZGCqINHtnfEiAns8WXlA8t3lt66/ItadIoPG6
dQTgqepcBKqQ4mUiS5UKPO5GTGEe43ZWTR8slXX1yd8XwiUL0PqTu1FDERsJbm/1rT0ehNJOBpd7
zmtnv/nJDgpuIpDKG9LPUoB92VW084IgRaupRcylWyxLXmCYvaREVljor9v5l+hZcQT2d5B5rwO5
n4ukyE2hSAcs6WUSwy0AMB42OewijayrSQ5ijprtTfrK7Efei75qLQbHBcDaXWWTZ/hDknebRWsY
IMjtXtfA17rqu+3BfB+T0h+zMs+IEfWC979yHZAUhT4g4TQeOuOVZkfKmiclP28nPWbE3ox6nNEX
0B3DpWtRBaMrGLMwARCe0LOnR3VoaP4A2jKik6jkSfZQDDU3IdNd8myd+5pF/qFuo3KM9YWUhs57
f9skEVXtmreeV/LZQIi/U9a7/jLdJVaN5x1n+MSJkicpibGSfGaku7c7nUXJzVDQLVxjn/LD1JdK
wMCD1Kgs+7/QnyYNtRQ+5S7SohzAm9KtUUYy7ddjI6So4eiulwH5wDeNioltGk1b5nJkVlRavKAH
nNK7w1CI3loUOh7EGcLXNlPVO0SS6oneGSj23Zx9OmbD1VABnVKE58lSJGnD6J7G4PTfVJvfTnr9
+1ZFW/IVQEO3LWSBH0+iUc9cGKVS9o0XjemlN27AyvFDkpWElz789imCl7g+647KVMxLYqiJdNrw
XnHKBCbVmQ+v0Wwi6HkUXmerAWyVqtDnioSPHwFOrZzqcjgkGsi0dmm7bkSJMkeJ4FQP7RtToFCW
eE+foZLCptye3TSCSNfCliVyCE8/n8MljNJW+nHdRx9/hVVI0Bdt1gqBIoTnhJrSfp+lBasj3RTR
DBCJJeEFt4vw0fOI7bvlgqfd1iQYlwkARK8KH8PV0cjSmrZn4i/vIZJQE9nNNu2NNwcOTMMLERiC
AaizFtlYC2HdgifzkPUre3JWLraeoPM8vWKwMXAink7X8N1tThh+2hJnRSU9okyTbxPV9AaeWkX7
U83jMLDqy31MFeCes2+WsBzpeInfr4aQ5do1jnQzCyAbAu2Bc4phxEhFB1BmMhrJcIJ8YoKyMbRk
112ZUSKnBZToDn/b8xWPNs1+j7ovfLknKktcnOPk5V3Z97Ro8MTbmd0C3xKR6+QxDVJ98mOl8x29
Yhr+ej6fX0myY7y/arcjE9f0/WV9qNXba9WDkGB+Iphrqf7uo5YL1QaYgVS/1kBVUBY+OdBPnxoN
Ns7KyTG7VMj+mdJx/d3NJZRozs6USBHk5Cj7KUjRhU6/2KZeoRlZ29IPrBqCxIVdXGfJTrjCwPzB
icD4EFGani6RNj1+gN7Gpv9NmtNWeI/edEjb78BOI2GbXFvq+0HNvyRZttSYW9m5TNc0jcHVOTQc
EF6jebNY0JMMHyLQRohAi01Qtqw3S9cu1zSVSzQdANIw//K2PUQP0ShoplPP7CJOufxDiCHV35dY
O3qBB/5/nXnn5ZJ3N9ev7tg+2+km3L03lqzPeldRslPNk4j5ldxKGmLaYf6pLRWx2SqHuDJi2GMd
09AorQguENQwqgA+GXaWRt6f66CqgBV77/W6kUPifkoFeWgphsOUQLrAgIcRjIc+gJ9ZFOMBaanm
i1CkasJq18JEeFNLasgwwZKDI6R1mwO8GZi3LKGKCxIXFQIMmPsi7TsX6sF3W0q4IyaPBKzjwXIP
4UY5VuinGCPAXwFgq+SCFLJDh7aG2VWayd+nqG2J55WfLhe1nj3vfApFlOTISzEa/M3oTsMovZ/T
KzyZXt8/8MionyvTp5s7uX/jEgaDMQdcgdSUr3h5a/SOb4tG7iiOue7AwzAo5xKEyikQ3XT6zBi/
n5GadwXz8iFVhzifdgNdvvv07tl2A35gKBB94oYr3y6R5CFqJYleJo+nzEO0XrtmOcG8n+0Ropnn
9yMb/+K3pkcfWlhMIxBIz39RWZOzSAOXhTJnwb1n+6n1Yww3ZK3jZtmzpBEK8AvYg54H3wG45YEs
LFzyFVLykCtBGYGW6xPPGaJRVeBU/O0+9MUcGxE0OL1fiPd6Y1UELof1TCfylBYVWTujKxJetRW6
YFmDNl63YEA0jpx1bVqw0O0lBhe5dZJl/9SY+pTx80OOpK+eO7ghjdr614rotRmB8a2dlKxqYUIs
a8BC3tonesB5pPsUIMQlhEGg+IaZYbiCo/8LMunXaIoxpyxoyysUlZ6vChOZtLaSoJ4KDlMfxlJn
/twGFjyt2VVuhZYddI3Az+gnoLZZmhisxrv6u65jDA2+EyT6qkWYqVYZwygCK4Rn48YKtou0bapM
0V/28ZBUFg40tBZ6CqlWb1FrRRWuxZdc63GDmidgbBRzFPr3tog6QdDi+PuS8etS7+ofN04HiJfH
JqbqnUsaWiiWV2VnZSRTkZsU9yt+1A+hCmoombFsUwosTIcx6VavNSJs7rNGCNrN44czu5PoR59P
ki+HgjGu1/zNIpyB1KgKK6slldBlG4olUfJw8PEi+ma7hz8EGzxsHH/udxZ/yVOX6p++OARbdMaz
ig/ZlyGPQwy25x+0r3JH01qt5bxM1WWeQ0qVyMOwSBRBipos4GiajgZp6cnQKBCFldRA3fJZlnpw
8pxp978onOPDgpUx1lWWD3NdVj12MxUrxALtiWDOvDDU0fzpwGlylARf+mexzcjDwhV1oh45rZAI
l05enW2ge7GwZ3CZdoRFo5ptPl2MGIO6flCEfkafXMsutyBctsMfaYUl9oRtHVG66XlaL8oIZzXZ
6ZxfBJJWWYgFyES9/7Okpnyn/7M/LiI3Lo5HtlQuFj0X1Z4vF6+xKFl1WbKFB/b5K8JiaYODMsgA
RD3HZ0d8mZ2sdUV2f4053stgbJrIMoTsnrhlo3NeqwTDw/inb6MW2aK1ezz0QkzCEnE8qeKEcBU3
nEar5aYQZpZJcJZ7SoMBgJBfGFf8OSXrBJdFJzHTWv74O1Jbcd75rc/YaZGmu1PC6TG8xvlEm7z8
0QmjOIkkLZ4hE0Z0OiFKKMhIBhp6yUuEsdS5rC8ElFKEeoXgRep3op1BgPL7BKnAD9vCAUGr/2vc
c+iJThnzpDpzh+g7gcobTCq0QvXoslqliDY63uTJhHIYPVR5mLCEoAb94xPldWcPaMqNeFycx6Ky
oQsJ49CGkXAm4ST59863ESiT8aYwYgN/a0NfwSRUcmpoteUTtW1sAoJVU1D/SreI7SyShsF09GsD
5X9OrVQaonEKK3YTV9UYApOYBaSo9sEaDanynULWjo6NTNvB4tQGh4qN/2aN7Bxf7HBkMsZ1FnTo
KnqZmZ8+30hKgQ/dh0cC388FwiGGcM5o0Pa8/VwPRU8lpip0Gralx7gUPtQ82P8ioq3soxgvWNa9
yfmUHkdmUgJyaw5nkMOGmtqOX3hD+r5eZ6KWGXM+2qogj8tZDSlMLsAyKkZpT3nowg4PhxD2/Bql
oz5kqnQCn5pXHIj4Ah1pDSUNJEE5nkeuL9LKBgdtk4kUHCAqAVGZC2r1ZGj5M5dc5jEU9GCI5lTg
6izUraWqrwRguhmnZhCDadcjNYfdeZsrwuSVfA/HUAE9XSv9haPdNFWEhNgSdqMh9mUfbT+ddMN5
eTF/RURwKO19qaquKnYtNXYwOZaOjfU8rSjYHdyBalnBZ7aSM5urTeIpupZnM5iSRtfMG9N001UX
p94tfFGgUw4cDU6bHgEoN+5XUcwuwXC6oJCzAjmuxkIjHBjSdbYE+HeENy+0GAkl7Cx6p9nnMdBv
az2FkS0qCFIGxRDL3E4H28I4dWzDXqFggfxuVzE6mfO8adBW2lux0mWPft0XD6lKYwHu8ZRKjYUV
Uv4y2vid8Vix47ubiWgdWsTnNlWvGE6W3xOOjFjtby+FiWuvnLwMzuKCRITEcsAZZ42Hsvxvd+HE
MHc8M4j/S3OeHYEl0PSFq8QullFwcZYKdVFdFWJcAzX/05JVBEWn4a4GDCgMEjTuIzC12+EsovN+
ZG9u6nNuNuNV7w91tjovRhqF1fvMKLy2+cVuJmlTk87PjnyWMlEuxj5rQWWa3BfMMY0FZTlNTn8L
hvizfs9E/1Kp4twhSXC69HE22Tf/aoWkAFTnD8KtuUHD4K2pmQyYKA2DabzBcEDIfJlQE2iaJVKu
PulC66Q5joX1prZNOVk3YW2egf5FV/8xdQVMK/4Cy4BqC1f2iJcio9kBloAcADmUPz1DfjQSoh0k
y82AovkhLuVxaGu1Il9KqH9QM4CGFcH1NQSEOEvA5kjoAznEeVQUk/D7GSPxMr4xZqVtPm60zoYG
LMt+xnUGn+L8kBU3V8kIUkTXcUDJ/KwtIv3bGUhSDDjJ24wTCZXWXjHCAzB6ofjfaUF4bvVuefUr
P5RCPfAlyhfI+LOnR0FCZVHpZBUxgmDVRW+wt/Y4QvH8e6Cz1k25Q6J4/YjMkd5KOiNtRSbkVds5
strTqTn6eb8DG8RvtBMkNuxtCHKyhs2jVsHTSkc2UjOxHYPN1A5Rpv/DMApwUlo11KcuBfwnK+fU
admTz0aE8s2sdGjcTezekpboJLyB2+F9FE/qZj/IutDcHrefgUqhi+MfA6tcEsyb7kX6fcdLZ1zu
EBkyo5Z+PSsRaLG8/LLQ2NDvAEtSv1X2jIB9mw8RHVISPcQN8xliE0IpzQHc+UlmIqfmr/w9gNQv
IFqIpDJ0eGUEIsn1sZZfvqJuuL4CpJoUQUe/x+L4jlfnnEMXS3kqiIr445EFL5WwavTF6Ok3rT+p
284twpa/b5Pdm48OdhpNSzLtL8jmFERkkpH6C4i4M5U4tjcxCE1ITkQYE4OUe4io0C5uH9tuk9uS
CYwgcd0iB7X2AeZ6m8Py1qwtipozp6wgwIV6Wy8WtIrFYehEnlR1KSU9+KM1kEk1emb1LnnQsHxc
pe5LGybYVc2LfaY2xkcwrXR885dklhdvLoAy870EzRS4JNZwr+w2mT+Zklb0zaM8EVZPKbhPd9xC
v8LehIEqAJRyjHgvz0v9jkS+X5o+OKNYhSKgG+wT1IuMDABFObbCLACmpvBUMZpjXrIL9a0vNgDm
GNv6yQnVSJbsQx0VFxCZuhN5el8iPqS48hAMV+fZPw3Z/is9hxCcbko5MnvdyMs8oPF/xdb/wIZe
MgQAgWJSYdLxLraPJPN7zrND1l8nIkcBh+7AcPLXtYXI9jRsVzwjFvn9UkMrtTnnMop6IWW6Q4nZ
NA8B0ePBa+rON4QliTlzT/wgd2gM2IygXK9qxlOVjsq1/D3nM3MdE7rTWVOVwRStt6OBHSnlXJr4
MlDapLzYQ7/bfN1lbOap5fUoc6nRPLzmsN42Uhs6/UHuDvB+zyolbIPOjm+eleLIhmrPRhbDojD6
e9koi/AxwqFqIeUiXWYmFUTHzeiBdeWse/W/iiBEVXyNopCiFYwox3XOedAlbQ3ZgPDEJ5DtiFAm
koMPAU5Osxalt7vQNnd0crUiX83lDVNpIo6AJWiMjjLh+KxJLoNl7aLQGB3SKTKjC0aOdHWI/V/q
j9bDU9dLWI8VbXcZz4r72eRC7ETmbzHw1C33y0+fCErwWRyBkFLZW2yMN3ZryMy4depVL2de+6o5
AfTJbqgJsKIgy0tIQ4ae+UTwpMzRLmBjOav/LP9FIdILKSO+uYswD6HutYZ9x3o8RAjyGGEt4QGQ
+0ilAG8FxRUF1RZ2YBXQdZyi5WZbSTHUaQXCWfN2FVYPJXGOV62QZV2v+s5o+EpeAF8Ewi8odGQ7
3eclKwyRaqSJqrVgWUGjhg/YtnRW94q2D0ZYUWPrivTcEENmS/LmcY4X8wFkcjPDnK1dDUP0u3N6
4PaMKRPEgxnvMZJ12eLBRaZEgjf5A27NtY6AdxxTygT1KiZMQhOK+9584gE5pNKvtTP0kvDeEVm9
3zzFhtuy1V2E08gCroLTd0GiWg1Uv/QUkuy03FAFT88h7LzUFlP4VJrYLpP4yWrMiJGqp4mBKqqK
zgoTBG3n4fQuIQC4jynTuvAXWOhehC96n8ekSLnO8jp5ZaIYq4p3S5Hx5HLhNSDRmUcVLKGrM7YS
TseOOrxvA0ghUVIfVbZUty6LtL1W2ZxWv062w183Ivbhwv9VPOT0xeu60kNaDZN1ukyEdrB7KflK
mX+Vx7M6Lcm3yVercX7MAqm+dF3ICpNSC56aMJYw3f9tts/mYBCa1VeFdPe3YiMRRIMxihJi2V9K
8JlY4FYit/F3UYoM4TWZwt3NEj7RbIJqmP21bNwIFqYeryXdS4ToBlc0gYPFVU/ehMS3eWzf/LMJ
phRYD9cV7hGNUluhadICQOuWbA7hqx8o8uby3ApSSyZes/QB+uYFND35Kq7aEYxzmDTVQPFQbBRS
1Lk2Zvqag3aCnjFPdgSpfMioOPyJRP1psxMhJgOToo2d3wXIFSZu5Jq+X3pIVRHApyIRRCfwy32E
x8hqQWhmBbIqIERYbkfCzouNanf4jKtn98d3/RqYsTaV9VeDV1LzsUHeRG4HKH7SvkI+pX/lj9Nr
Ex3ugw7Ubh60Hq5X/LkTjJWpSVTzqHZ6r3NBMOmOhtjbVC9Og+R2Wwx9fuJHe4px4pIGAHYP8Mff
hj8DFIq6Grs1KGvZctOmVu1ercBBuDabATtjPkbx7jYuix3eIiAfErqaYcHknL3NF6Nij/i/3PWH
4rP0IlehQjNJTwBg/bY+9HPdimZR98ZpCNvnax0xHgBeCe/+sXu8Mxl8xnzB8npmS4SWBT5wC/ZZ
ed4Rv1m7qBlOWBWiSgfCANtYye/amP7Qm0u54d2RlQ50uIXAh1XEROtVbq0aANrZ2z1QDQOhNMi4
TItz3U/gGaOr5yCLta/Q0jRzZaLjaFsw3cl8XOaHmZpgOp31sY2aE61lxOnuKTDFRkHfqRFMNYCT
oB9q9COBF7TZxU++OiXhI0uf0RYHR2NphgPmFkuKkvSIK+vW5gzQp1hdBk0m2vZPWl1qywmWe5V3
UhSD2wyNUHjZsFY8E6Jl22R7HENmko5ESdt+A6C9QSdjmqOJhlmAAyHYr66jcQCeD/DW3KaG0LUy
9lhqS6hGNZJXTUbVGWbNt30cRRUXLXHtmlKYZu7QhXNDxE3zdd9woWRCkkhBDoFpTN2m4vl7ERIx
feMBcMeqxh1dqqP+RBZ4klxWhnIl+D7BCIq/hEVkkinsUOy2aklwugOZI6jdt347UsGiNlwacEy2
TiCe/f80q7SAT+UheTNFJuZJsani+OWp0WF0b+cElVFTMyMcro5swnpbR3fcXjSbOmu7W8yDU564
wRH8T4GkbDpRd8MOWxQvb4yw4HJhly6oJQMypTK//w+n9vdWyvrvQbgHhqRZpCfOwrpdMnGr/M0n
GwQdQ59wFeubFSU7k9USNLmkame3Qnq/fR4U7CaZGc+L/TccvQgpnrwQstD3JTFMA3q7Vi/C1BwE
pBxST1lgxDJEuswEzklhKr/e+tqd1IAH7v5NcrvJRzzq5kYkVHcz8FK1dyUi3SgUbp2CLCL5/rV9
kIIgeqIgk+fvILAG1MrYv+sfYuy3CXHFgtNMgg63iV4YqbBazp5tGzI8mF3Z6IfNrFHOwqJYSkzE
W0Lx+jOrjWBGHXKXT5Jxw6SSBWtBjorPs3ciyxM9omaNBO6gYsx5/sSZJbHj7jujMhVQd/Gr08+C
S877H5p/H2xGEVwnswXxcFOYMZwp8UHY5/X9yL8t42ekAOlZNr5WWNMxWQjSWpiqMqnnOSG+bv1H
mRFF0hVig893RmyQgWxxN2XlO99L/bPzeRIuWukNwViYKKe5ZVxyfD/qfMGwLPQCPpnxXBpuSmfn
o+XzkADs/hPSVqO0CrHaXyUK+arp2Lppgzs5EzprOUZBg0ou83sNBnQ4hJaS7J0wMUAj3LZt/T9o
wMi8Q1xplQVDIbDZkIRpOvTKfGeWQ5nf1LI9P4Wk/3XDkMDvNWyM4WNE+p1yvdHUSjHwk36a+AwI
xH3T+MEYyOeYkinIiAN6YrAhmYtqYMGqYOfva67Np4kBe+gf9tKb9+5/TKxGFwbS5sFtGbLNCKkT
ebYVVgPQpKQyGBVEmUr485rMng8u6HzocLNa2v/mlNnlw4aS2asAHBAGi9ne7wXWePnTFd1SJHA2
CrX2x1kefgihHa+rIdKgRHsMBbYYjfcHEV1DBIvVGzYDM/OQTZIeKJOpjUaCe/7Id/EO8Ab94de9
e1y7mX8tXNw6XMVZiXTTczfUZvFNJnGASslOVk2ynRqzCfGjCA21b23ylks+p1OlPhyzI5gOxeuS
wo02x9h7iK6NX7lVyvCpr2dVyXt6TaoAce0gELrQE9CxPqB8D6LxAZOIWFaQYLxWQjLM93TgjYY2
3V/oGJch7XY3t7UrzUyc/LXo3dT4q140v6j4fiEV+i+mfOEXTTSzmotCb5AurGzWPxh4vANfh4dj
n6JMCuom2A8oEcxTXw7zluSz0To05/p61E6V0BhxhEdiBBU/4UiVFPN1Mc+RoPkCkVUcnlahj8E1
chSauZ/HLRtqwtuCKLXTW4OoSCQDA5liQMOcyvdd0cM8+SCE1vKrkxch4IlEFqqLOfN5Ou9pFT2B
plDxGmQeO5z4KuEwiNUtxRTKXftszOnz4gnIuUlds9U0XCIYE6+5bCvjpHXnGCdgJ/urlqurcXnG
zcA4ghbje8b2gomBq4j/5sH24ZAGlqOtW7qqvIxk0q/yXncPrbHt2ERNG6nVtWL+yxv0fMRK3d+l
iAll4IA+zIV8lvMfpEgwSS+3J1NbwmyjKuSN4WO4m+IkRkGwuv5LhPVs2SpyUlziFwjcGEoey9fr
QTQC/IpomRgkET5+cAHBJuNJ4Wf0IchXVJ7O+VCwKhes7Q5DnnhgyHd0rsxt63l9T/AsJvJR5on+
bf3rZNjCVIKdweJW/le9iRKK5IuTUm/73fc2tQwNS6abgtEviMsQw3faHVhQaf13PyARMvAmaKg9
gTAhM7efLLgb3c0yoAJH4LMP9vSp6KcPBQAs4rhT90A85T6d+lLRQYOu0bFVgupeuWs0C1ZFzyPA
T1i6TRVx9rrcrtOZ15Dkck1XJknfDpo4Usa9WyBlDiFfQISC+gHVaT5ALuB471RML9xY71HuWSa2
SAoWkFVOuZjLAziuJpRoGP6u7lDBRlFUvp5dk7+yGpm/4xJenCt9hOCiMaKgkEvp6uy3ORrRPIEE
nXkmYe3bdcD1iZVov5u+Yh1TB6ASB1qmsd6LvZ2doocesUFRzrDBQMGFiDaGCdWPbAftdvJJy+3q
8iZjKicO9UEetF0OydWQZQCkGBFQ3eT5jPdOW1K5aCxciNUR0BvwvT7OsiAZixNg+5Ve7C0o0Wtd
SEHD5JfQmzkSulLjrSGOJmLRgegOtqrlW+2f6h+a2KdqQ1/rQTyW4RlCVNoFv47r+7TPM5RILaSa
pnqKC4lfFZJuzNXd8CI683EJIorc6AL47l0Q++i6UdI/tMMww5AJrGyzroKcflu+aHD7Pt3Xj3Tw
fEeTku6ElKl1QgS/DDuXaKhpJkrwcQzYtGYMd8DRetfAU/sPwEXLdLlOKGmRi41ZNTA3wofKqUjG
xirmKxhzk4CsWcSR+5H89SMDMx7zAcZXjAoGjc+uQYiT7E1bGJ6rzOOvZ6jzJRLEig/nJ1wj0732
Utsqnrv1UQwRqb0GkQATHRhAWOYd2A+Twi4C0IfHyY/OGKGhxYFey05b2VJmJ0E56pXfn1PCRwoC
CoUUxXH7a7KL5pFtrlnc+aMznQ9pEK97rv8czr9j60vDxKc/5PkQC68vUFkfN3szDr8J3GXP2xlQ
hi4jqOYwb+AiyUqQBxK3FKSC2qa0OBLEgMebLTlmVkhFvhiXP02q0BMSYILNBiT3QKAkAg8gJ/YJ
GCbtdpa+BMh0LfOKiDc2sNVEHLAUzjQtXgn5TFPDNvq8tFMjQAfqs4GPiubuejn0zbHnWhNhMUI7
19NXVNM2Fl9+JpsA3rv233UqnXMgU5+/rtLO1wkUVMKWvu3+iUcLFiYNyDHXd0lUAmUw3aSd13aE
isvJZ7A1EUHZ8sGspOqyfxWM7NzdF8F/jSYpl0hHw5xkCLtrS6cPQG4NtgQs6kXCf40ExLQ2f0R7
n0I44MzcusOr5/H9kANWVAm6Q1Nr0K7kKnoQP4cU9T/pJoc4SaZV+J9bOa8UTbZPzrcfZRp8s4x2
CbxmGPbwO3Nkkx8zp9+pINkwLFVsPHL6DHwGZtmSAqXMyzw/2uYJzJlcG9dfq8yrEtLQPR//Hqi3
yB+L+eCL8Ikchlda6f+rjy+qQIOpcKQLzLste5KeTxb67EMWcauV/o2RM6jkO6nrnayuiWwVCEgr
srNntT43X47mYowfilsBwe+tbZKf01NyGzSQKJt8TxnNSSsRmOzaT0mzEyZA7Ug5AAC2h+gvq3Ds
hQe3QK3BWPM6vJki7HUz+Vtdww4MrGB1gn4NuRbeW+d1RqXeDHx5T9IvKQbTJoWldNmw2cbGSmaz
CTGtFluV5IbS9Ym92BcmYn07r2UFtyECRKiumaGVNBMUYdpbVDiDua2yV4VV1VX9Ya5HkP7MS9o+
dmKxGvt1FunfXFEYAcUNiHr/5qdwjwOFsoKQd97Z8KsMTCYbS5lNa5E7I2SEUpf8Vro/VT+FNx+Y
8B499wWLxvdxult5TI4J5klpTm6gYu9c/aBFEgaU7+10wakEk+UL1HfzyRAiTMAVu6OiZSk0nHEc
a6fwMQLp/KSs4zRn/xxloyLrUxTZk2++L+E0OU7f3dFCXt29UY9+aYg4ZIh2BsEBJob/0oS6G7TX
/fRDVK+0zplQxP47mek2+S/v5EmQAPjGPvs6k68vYGQ2bwqlhlH2//ttyrBus+h8vfjYjRcBOneR
mf0GNDakKkmalFlNr7XaJeGUMVORZOAyBMHCB5S5ccCYgeMbFgbV8rx1fStNVH1a6nVDoueHNI2X
YI6maF71zyTZjhM93APxvM9npzeu8eoAejn3eeQvJAju/50n03Bi6B9OoFYZZOCEqcaQgnOnwdHa
9V+gG+BHriW0iKDBLG+ZLnExyOG7Wxf5JBR5JiyeX+k1A24Ib1HKbQyuXCbHPAm5HUjul0NcBooS
Ps5Q5RnwEoPaD4fH2I9dt089NZugMqSrtemD5QmQRrxPhLWBx90z//GWNwLL4z8zClKAde2KSWPo
/kV80xXzaIvyG7XnMnlYsMaPyf+at4KMV975sJqk0dqNmQe+d0pIPoz78MCR/9S8dpS060/A2jp+
LIW859HQNFGRl/pmHDq9dwiQZsisyVRTFyZoVMsRmfSUyryWxG/p50AxGceUaAT16tL8kQAUbe4x
a02ulKerSt+cA+pSrnQ3NmDxiGkPMIDZMVuR+rNHwcHpuI7kbDre/1k36ju9qv1iu8vMmz257mIO
l0hnyrCblfRk1aRa2wKxY0XU+wrTN9gFEF+DD5iRXH3QZavZtziGDi7uDCpwek16+uVOPyFNMwbg
nN1Na4UU0fJD26ZKHG7dhdOd3ZWOtHjWbrQYcwZJ5Xv3TdkHSjjKLxipyH8ith6nXl/zfO46Oo6Z
SrR/dp7xcgwSu++MtdK6ZswSjgQyOHCIZk/L/2Z28rzu34o8z4HBMAkEpi6lhQXVTTbhJWfW9pDZ
PtUIatTNJKQL1F4ftxp9VCF7aGfrwNj1BtEKHgvZL15FftXjYhEDuA3cTgX9wDr/6tV+fMFDdefI
ak+C4dVShgbYMtQ4xOx8MfpzLzmUQae9RiH2D2/RZ+o8Qv2a6T1rIOl2a45REw1pn6bBOJDOr+GC
DyOS4FyEFZD/8G2adzdt+MSju7CK+FQ2W7iq9mLtqud/BuPyn74E8GB02vZduM7EfpNhf0mZbWK5
qSwv1fUx+i8WPtVH/p7GEWL223FJqP3JuqJYb/zfqLCS5Jw8JCZcykpU3n5nTdEOM0pGVgXaZIKc
UAsNn0XqhEofww/VYY99V+1boWH2bg4VE9nLKjcwGiuG27/Q9grBvF/GOqbKm8lGBbb2pJf3OIgZ
h3xe0q83YoYBYNkY5w35ckX3jlxmTu1GY9c+VQWHm25yBIqTOpiylU0M0rSjkXlG1KJxWhV0PuyO
Qg5Gollrw6Xewi0IYdb4ZdKjEfmoORGSETG5Aobf9iFnsQel97oNgoJO4eCh5Kxru8UqT28G6whO
1kbWWFJ1WTvJiptowbZnGfYTrKgBapYR/ncqjkLAXvRA6vXBeLR0I3H/xDolHuwh/MR9iiROiKgs
ZPnNTmClO1i6ULUgRQ/AvfjNdhQ+EdEZYmj/kj9DvqatEfqfBy2u/Wpgni1YkUO9dQY5CORcGS9M
tNYdIUlHlxjPA9pIB1XYTbXC84Pqn/HTkq5C8KJ73Non3fi3UjNsGnjbn+2nNdUSwSuVdqHGLfeL
zW3Mz1OLDVyKcennuItCK2YTA24XWvvUEDNVqFPCMBrwgOFSymUou1GQ9dC+yvRBB7hL9iMEczjp
+s/pBgMgwrBCZ5VYCp6NvE3L03kXTCnDdx9q8N08aTnDsMySQZZk2uGIKyETsI8dXMkdyzwn+TmI
CVpPDRvcLFw5HPksSQiKiyT0+jc1Twkux+ojz8BQDjpwB2DQEEzUwtkO0StpVHsOOWRRkLIarKxt
IjMLZwguKynC48Y+FaXjT6iAj1EkVGIVSOstbcrJ6V8uNBdUDCE4lUDDjQiwhVxB8z+/zT2YG4Ty
u/oOEMN72qWUTtbBctS2/IPLixB6OoksY3niklDUVdNEcpvOEZnwdiWK1oJXaYFhzc0DUVBZNp14
kHIKM5i9ZSW+4I1mIV6Mno4Op9h9HituI7owRexQcXElofbc5pKzrceOVSrZ7GlpHSbECB1Gm8yL
xBBAvad3VNUBlj4WzDS13jiJica9Pgc/PZEE44HsVSFugcedolH7wNBKP2U+NOzLBZ9GCsmHUo7C
qmNDi8K0jb4TDbPfwjhjqx+yf9cVvdfOaStgxhXQ2Qvl1X+hunInAe7IML+lyi1jGohiB8Qc0AGn
yuuUDWPglAy5ucBt9k15m6klmUk2OJ55qf3kUGnvixkACcx6AvnOwg7ueHDURvp3RnORRtgpO22+
HgTA1uTsjkON9ab+OeS5J2vdDqEhSJTrOgGyNWzZXAjec2wm2Z9GGQwz6FoxW+hZaZblsmYHTInL
nVKRUaD0452iFJrB4rD+BFIGyTjMJRq1jI2WhWOTIIOUw3gs5Zn9YQYwSlaQZhCqvFxiaPomCdb0
z93L6T/1oolxVvIzaeMWnCbGs0vrNy4w/hgvVbR1HvOytJ3YllOi9FKelKx05lgHUx0I0bKqTybO
8gHrpJRSTEvCi3VFK1aiW0FB2qB92dnkdxx9m4I0caLtFzYsizz5WwXCNdsPUVsc9C5zIyioT7AW
ustx8wHA8PjR4ue/ti4jx0vNDoanajGS5YzcIPzoOiGeIjGJzwT52/91ONBsRJiYOZpQUNaKPk2q
JGnRiR1jhwETgqrXBOqaaTDPxtQmlGDtt30dMe94CXkr0Jqy+8YN7OLWCXavtsZ3SY4P+QRZf8CP
LV22lfFjQpSX8gYIF2kVKZj0szYu5jYka/56BBi4DHZ2AU9o8/ofR0j12NRzUiyhvJiYXn2pyEB3
BvYMuzEHtIOsVQi8B5jT2M5FYtsxQWC/VhMPj759io8mChgq4KiJx/5JtZ5UvhxwFbMrCxFnO/+i
7RR2HzpGd+WLjWmecNRF/U4MrF32sDHg3T7vmSK8wN5GYpIZAWexfVGeoVmRAIlCWfQqL+h/MVpH
1OwuOnpsqv9U4LYnmvNupmarhbpWwsSwPIvW5OKAJ8zhLBls1KpzoTp9CdFmo6rdJqDBfUjkmeXz
O2wkg3/R5wqp/J8RXXuMADc5BTSyzK6WRW77wjCvr2+wuMoZBwLJ+ckgHJM41lUYbwTuSQkEhHN+
u/B59mT8wdFL1nfRh2umHPVB36BZwWHyiSoPNMUpn43Ja5IVnaTAOqJtDMs4eL/+LkeD685jsKuE
CxuQCHYToYf5HCPUYLr6+fg80RpZUPWymH+DawkxbIRSAd3bVHhEvbTm+oSmFeUduulUczOWwyN7
xSlkJ1oQFosUf/2ceCiZ2ErPX4PWegYgBi4qYec5mrZL0Dc55XGCKLoEvnSVE+PpsU5mXfTTxKBo
COJ7NBFMoyEHIpShTu9TApEtnr+n8RO2g7SeUK04aVkTj9LAt4zUquX7lXwuDipJ5O/AQaYcGtlq
GY4w7jFFqrBsYAQTAbIm7j5bNlPWU/OLRqx8jNG7QA8hCrUUDHhcSSrNFOqP8RGfiBuSMkFigMIo
8Cl3lNlkEs90MUxT/VDUNWgrClq92+t3Zr051X8ReegWyeGAHKYfNGU0eF/yu4UIWacCpdpzTJoQ
sSJGWwITDy6M2//BqFkyf34gWh1/uI23oN+1eb08BPqNqF819xlqsYP2kqhu+YD2zhl2FgIKptDa
E5+KwxJTA9u8HFH82XM4oi25ZdXTax0P5zEBEZql2N0Sr6YksVycGx2CIvQntKVYU/3IPY902bPm
u3YS17A6+M0BRaICjuw6LYct0FJDwqfrskpAelyXoJQZdJOTtzUDwKvPLXqgBZtS+hmwyXvQ7ziL
jXfGaqhH4EoCCnymb/MMJSBzRk+tQMPnVki03Pk7po4yimomNlqsy+XZrBZ51L4yux0hRnvyfFsc
/o0iIVTSGYPl0O8AU3VfQbB9chjeoCczEkXKNmA2HYssi8LhrcZ7H0mDjG4t97fVh1P11Q2TbMKP
LZIo2PmkDO1++b2CpR7hMjVEOphjb6itK8YWkjsQf5OT2pbOkwXv0y+Y3Mdj5mm0tFhg1P51nIsl
BzBj/kxnGS953GbjElQsYv6WSBoPNkxMxlRbBFVZXTX/vYapE8L+cmpZyO0TxjxC3LERkTUWQviM
bnxDHKEsdnU7+2ykcVD+fPVqLYcHItxbO9BrgVSLQTEAoArZlL+ltBn1tzriwJ79TyILL8xflvD3
O5y9QnOkwZ31NZw/rw9HNGkkrPJXuqfacbd0nEZ8bB67bCwemf3XHLfryO9IYnL/gzRZht+It8bK
PvnBRwvAIv29n1a96nmMrEYuitvZ0gtBoLQxI1QtfqGjwqJq2iFmv2yaQm/S4W3kMuJst4iJrWRl
wLNTe7GCNHMaYwEmKNxvNI1+hWYFAHAx9FuCDulbX4wTBrDlBLeEjzzK5Fhp6CDggbRAeTZEdpCG
VuncYQnsszHwT/euTOkCRCCg32zRs5sNOHPwExDrwgU8wBCZzOvtqz24CnTXBeuVDTJuEWpqU4tU
0nSNC7eAztbsSXzl4GIuOLfWjjhCqYO5poKEoeeOmfyFoiWE5GxlGSRVPOMuJ+UZjMgJqWxI0CeZ
qaP5eZ3HQ0PywRnP3HkZl8hUV684aSR/ZpPw3oF9Z0TDzSu2uuc6thdZZkJAklVyuulhVfwUM8oy
nLKpsvmthnt0FZD6+PtI544as/9h6G0VEarqLrl1vBelhkURE6VJRc5bsi2ZbWnUhV4fu6VIy7e3
NIg3dgmnO1kdPiD2VTH1nh9uzl9gqSCvSQqUm9IuNyhz7xe5i2euF8LvdKiSoOlK1wuF2M9GWdE/
CNqGEEmJgWcQA9TFgPCv0RYQ8E+JblVskROLR8NaRGcy5MbAGk2KxHfZqSa50bN+qJuE73raOZcO
7TL54yHIl4OGnAMVG+Eaia92GdTDy9VkXTrLJvAgKcGiGzHaxqXMfcXW/683XvJWN7Ir9hKRx98W
TkEZnLJfiQW8g55VmbdMrOEMCbfJKaRQzo3TODoZW91fD1l7m4bILKFQ3OuCNyppILmcgpVqIjfK
B7dqFUuXXNbkrD9bC8boL1O2yiD/sAiduUieqtpLDGJmNpnP5j6TWmev990s95DyFtPHAwircmuI
GEPb5z8S8re1x1F3EQjvRRekvsFZ9plVpij/W7+kaYElZyRsFF4CINNhMD5aSTThfIRkKHgYoRz+
W9gQm6tSg4HarPFXKyPVG6BDTJAWT3TDL1wKtj1vOeru+YR9M2Zg49JHU3rxoRwXc23wHERKd7w/
LMDjw9V3lqQCdsNZR2BSjNOOznhdZvw5ZJTGBWcHdXwnLZl4CPRpjXRDWd1CE6Q6AlNvAE02qDFN
rPlf7iwNnkXX1/yQ42CuqmAGtJWJSTbeN/iCpDf7wq0OrKcb/PPMP3nRwvoODr4L+k8CrzJ+rcn8
4zm6HG78bD6a8fJi8jC+TeHIDCekCcQihzpm0GwlZCfw8Zy1HFwIt4urhEfm9Gl+4cw6xDG6obWZ
R1hhEilUGfjOYrAHJiTx1IKBAVZlut9uAjjXAASAiGEeKef+sfWZIlX8mN12dWE0XsJJAG2Dk5Hv
yfsvYNzPE5Ecl/OO4Oveu9wZPWfIje2pTHt7fXutqH9+HkFxodFyHuOL4LtH3qQd8fepZVx2lAT0
Q77fjX76s6+01XpEZ888PpRxrp+m3ZoC4VhkuMWR+7U3FSDdqpxiHHTfoxJ6sSlWFVXlc34+WmrB
qJz6+ALJSYxgqe6CFS/7xMual7ct57O31crHPUx9nGOIbWuZShpXdzFHKuo6THbbFSn70S3ZUOlR
CI5gcmUkUVM/k6U/Vf2KbceZO3urFFIC3u0tB9hh/x44cJRj7l9ccnI6yse+Gf9k+6I5xO4fdXQJ
5wzBoF0OHiCercpWIFeDG8BokVhF4pn3bsfpLKeabfSPOkYXkoJc5r9QGVO7I94PmMZg4qZAcZat
KWeUacn68oC7QbG8ODBQEAvGVsXJZgudCs7mEGo98DIbCM1OyjLMxfxIyldH6NBCmJ3nFmEMswHz
SfUzBX+3z05EjTNBqEy7RTNSqvg27HqAmn4mXyVyrZN21X8Kirjdp6XKaqnlIgk7OCxNyWh+8ko0
z57/YlNQXRNIOdKdKYUGcuxxV5063xrMQ3c9LLr4gZWeMJZ78/328FcThO4/r6A4iC3UNYKpZ6y6
DxEzf6DuIcusWtlqm6G2zaN+fPiK3pthTxSr4LnH60OOVe6U/1Xz7arZwfa+tDQOpOxBV3utt19J
cxtCx4Wb6OOoyrQoGQi+RRXGHHP3GbrUTiNed7wKyKKExw4Psblhsg8YHnSJ4v0nbbGILz3v4vuY
oWYLCX14ZEAyknSdDJOB3637PHDwXJ1vLp6+wTScHhUnIPvNcVQkRdI59ndPS2+fPqGxHKX3YxGk
547mY7pJSpmI818+0eRJiyRE/AeYD0+LSdWYjvfPPLK1Pv8r45Uktqa30vLa2hQiAyqNNb7D9Osj
LsDA1Bk2i4HJZMuE8WwxDy5S9jV1Ewg3peu42uSC2Veniq0RGputj1WlON6oTUS2uC2oTm9jK4c3
ckGm878mflOhzV2AuR0iGjag0XnXWLrSuSNOJjJjBGijgpsFiakITEkd6uRKKYhFat6iCFSrQxj+
Bnl1ZUMPsaiQaXa1QtE0R+E4I51lq/Y7PNESZ5VCQJF9xThiFHaKn9ZAb/JFUZw4L3SiIkvqn2Ye
Tc9C5gdJTO3b5C3E+76HyC57OrGMTotl4pff8xI+b/cuy7QRnSEjgsRHx9PRlucIbat3DNgmqDLM
YmoVihEJ5wH0zOK70VTTTnxBFZf7NsAa3VZ75vfaDsqxMoh/oyO07tOlmwIuENVKvxIi5B+QGQrQ
wKklqCijBdi5DPTDiNPuS7f6KWLqTc3R3Djdxcc5aIdb+E62bMwo2Q5Jlvb//AUQ94OjrlMWaRAI
HswEYeilIJ3GPq1Qo5wVJQc6UaQXxYGi/ztetUJekFYkEnFALRtes4sTh43qnNeJGRgGawCL+/h9
VDx3lfo1w7Rp63I16DYZVN3BQNFr4sNgwYif9o0NXfXTb2wVqhKEGQr1Ep1mpRCoRrykdyFEi7+Q
O6uaezlfQozTcERe/ToBFTfxN4OgoilRZaENiAwrLZ9RH0AKpqfpuQm8xTbV6edfg2nuQrjBKefe
BVjoesl2i8aS0D5cSQ6SuO+wkd8khk7xSU3+5RIUDy7nmUCeNXtMeSUC8+wUcEZOzEjK2tviTQ4T
Rn2HAc82LOkg7am5teG46Swj8CaUtyxBF3/nfapuWRqCgeEO/LkI9JMbO4cOvHQUo8B74LV9WqTV
NAWl27jzHW/hdEPi4/01dTgN44BrcRzoIPKf81WBSX20F8cAWTBmSNe1+HEnAUxGOZmqiOZGU6Ym
InBl/U/BkEC5WT3gY1vMIdvAMyyxzu8JfuvnSSFo9h/2I0WEW/tJtLhg9kxVRyzWrhhIBbxm1ghR
ryJIXuBF6e4ry9OZ+9zs/CMhFhwlBjdC/KmYtbVzvZB9K4KQskqMYZqT3un/O1wp687HDA4jTH6w
wirqzdsZRWuR0G7bUbbZaOa9AeMqpd+KXZdos7e4uuyeA6Wp5iLePQg8a5AJ6hePfNML4SAaNT6h
357KYM+DQsWm/doAQgT83S02TRnCxSaTRsBEw4a0fi9LXcs99UEr6BswNGcWZXv0GXfzpvTGoajx
S4IwGyXjrQgqSe2g0GN6ZYnsRWQSOcnbHnBPSFTKVOAaNRsiujL/cLq9NeUcX5ieO93uc+3dTCka
2hdD9YHrYeyObsAMFPrVCKm1ztqJ8vd+EIReYEXSa5wmBfKW7Rs+7HcOSphvIDQQ9J6MVV/gppel
ALuEsR3zZiJIREGwLbE4eUuK0t0uK5SrRdrp4wJ0cE9pC/Xf9X3lN1zwkZLcMwkMw5EnCqF3/Jy3
7AkNBP/FcW/KOp7D/ZcmaidjmEk1Ncxgq2udB9qsoSktEAz/W8xzx5hf9mKwkc9hrW4mQd+T5mVM
6YFSDqtAhlh9rdTP99ECaHuLFL3vHmUuJUj/H4y78ca2fel6b0V12ym+cQvcSDmtaBlfqtFR8yuH
jEGMp8rIEORySJxndxpXjJarJWl9bFrdx6ov4oWLgyhOluaWXtedsi7RB2maHYSFls7kR6tQX7Xt
bv7wYaFKQfLBXUB5lW6gk+NDqdN/zN5OfNSEBWWyNPf9VakDvsteZl6yi5uLsowz/P50ArA/1mc2
hHcY9KjXJ7pa88J/eJp+ks9uMPhOufynNfWQZGBYiOVhXvU73xKE3Rs2OYJ5f5UcAnYsauTSbboQ
c8iT9wa2Pcvf3EXn6hvSwgHQbKR3lAf1HV2EsRf0SlL+ZGQQ8u0eApeP2fBROMiM6TgJiMkdsUjf
8frmMuc9LmlpITcH01/sbzyj5CpmdT7I3p3NGCCkkVY/2SN9IzW6xj48PQdGY/+/LGLcTW7SP7/G
yVse3O0Qh2qTBORuUkk3WcktYOuSaayI5Qmxn8Sc8WzWKntJ4SBsOPMW07U5Fhk2B02mInlaiw+T
jnf8AGjqKy2NrX8p1TIrE0e5oJnccFnX44TLplolzHjSYUqgcgDLwqv/CvGWpoa0PlHgeV3XSxSt
HXrhbedcvnduMXZ2OAkBrJwNeAJRjM/ML+04+25APlaRKi0k352p9ZETfvjisFsz3HKnPNGmY63D
LhE+CKYAwOJVI5PXny1scwKh8on6lZI4CE4P/BTS6zqUgSzXSZBlPcK0s+R3V7pfRWqcurzDe5Qj
xlSO2FslysLbJt+LxcJp9GPdSmted/TUCJUoEN1awoy457ennrrGDchaXbEBcQR01OhnVqLBgMz3
3Z65+j2y9/pbVCC10FcmgSd49WJk475YZIpodu3//4IZm0/qviP+5hmjSaxC3sC2hKqr3OLAaTmE
e4USWJSTouHPOxoIpuSvKbnoxoMfFDqN8R8n5/3jdEPsOFLNfPLeQRiwin3wWWN5DzJnil7lf9Z2
MEonQe3qzCwfy14t9+XXaOWWnnqN+J9+C0ye/YRdSfQ6zcvDJRYuxDpCJJ8ns+ZC4g1xSTFtJIwC
rS95tjyXQg0n00xssxD4rBASvkG1KLkNeW34fsJeu/7rHkC7H7YDpZTG3kZ6+PDGCPjc7HqB93Lh
Z9Koy/Xrhq1rPNowiQfz22tEPRi3Hfv6dNzuzl2zAgVK6BRaZveY/LNqzOI4k0AK+NmjB4PdLUoU
LHX0+YuwR3Qm4nwGrTGash6SbK4dq6DYSpKtmBqGRImk834uc3bh2p0v6y+W+z2aUdunI6196E5Y
d/Ru5jcyYescqa9jxfzKax2CaQFYMNvej3dnoCnRO4vsxK/ZMId3qovOwo/OAE/NtMapQXQgZrRa
oYBRJFx5PXwl2Y6q0n3xmvZqL3yGmUOQqktLOU3uQ+h3vpmdF0S1PEbOX34L8afbGeAP8ySVmj0a
L6KTk1aTidU2UGi6TGaca72GW16+C5E74KGpyXvIAhDIUTkcMSftd8i+MqP5EKvbvtaUvmp3d33f
7fuS2wXjRLcmLE1m5Vg/noO2XaIPFMgtf43OvWSpvaQh13FLXgQW4NO1luwefKKiROKhze1/DTFl
IwLpcmn9UTJWap+DoHJgAMnXd289upbHr1prvqGpDKFYjcS4RYp381Yzpta0FRiRZ8nXrjt0U00l
Oe8VlcwmlhdvXkmTahQHFadYwL3FBjEqdCCpglk2VImKV95u4elfgTQp1mzfODqUmxw3dp6EzuS1
sQlsKt0r8eoFdpV5Vi4ClFYoAC26zMTPc2k7jK5pKoxL7l0rhS6yDrGbL/hrRAzbzSo1d9AfeTuZ
TOCWtWKHrcXOmzJPHQAkeXW8ek0TbSjDO5fe8yL35PrXRBEYOaap+CfTwhAQAIHhw4W5CAsJsw/9
/UbNamt5OZDgyAEzeC/numN/Szf8bApfeySHGh6v1A8ZybC3DT2jou8jlbDr/c+RqKF0YxV8nZ6T
A8Nuek4v4JB7lfhRv2jEXpVs9GU3/HNkHpylYfmbyoDax6CnaGbf3rxoxOqPJCdDm75WLalR+Q9N
HUQvxVxjL32wPrLGN6fhxlQcdoU8jcCxibYvc86pz7ksJRIv6P6Hl9aqeHoXnP32eDYXLshBI8pF
PQIHm1ZxwwAH7gkFSbYXRvffbwRaFjQEa16c21wtJe/cCMXKh+V95mLuZVNBpMSpUAczDSPBDwYp
M4T2L86tXnGT/4I5vI2bnU/HetXpfmq/IlPhfLbusxHay2C3YB0hR/NVu3e7so75AjogPrrUMPFB
cz+FoB7koWBLqAfOvllnl/2BBcD81HyG6nNg8QYEl5vI29GGNJ0yUMt96Iv5vuzA6HqzVPcp5O+G
j+FHhb08XGlNRxj4XR2FxOzwLtFKL83+7NkNBJt0IPC55XSlilIFaI885akBuaGNPJZvBFq+2FK4
K/4BqwoZARvxaTx3rqaqTEg/34lpMjwzfPZDvl8U/xin2Td3jhNJtzu654vNZ/zSf2FshM+mFhn0
bvxdr3b5vd/jr9vQzoGuHG5qOnO2AUzr3xf5MVZ1t70kbXtwuUjivlz/e3johzqAYb0qeht6S7Yk
KDqDSUz+n9fTyUihI3yBMT/Z6YaljVZNMK2cDLIovOELCHfnkYJRY7XlriSI77SH/3Oj3M9nq2NI
iCgD9hz/NeaaekX46vSCKH9u1S9JIRb2TQEYJhj9Zg/dsXc0zKvT9FKH9rGdiq3yg0z+HkyWKsy9
s9Q0vgDHVMzCdjlUUQ+hM/4GOnwpCK4y6AFnTxSPnodAGaKcuNIJq4ErlCOPQCkdT+7G5e0cqT/h
Pb1XRgszDbyXJN2ayHbum7uevgJy40EuISbBUM5uxCb9EMDU/SikzhmM2ICbq4aiQslKZwCZdieA
f9XTXebTvOQ+AMN+cZjDM3tFznng92VWKTpJp9Z8ULG3I1PmaWdlz6xvOfbA78MQvlpAJkac4MUm
a33bSCiiF1KLekziTRd2djs3EW1OoOdd80I8Th/8l07HhCcH6y1vmpG8RtBgb0b6xnnVcw3CuirM
rO/9Sf09TchamwymTtcLuzhFpUB85V9tt1K2nqondqAoRX5TWVbLkI26FPEqsgOs0Whcz84rIP3/
IjqpQaC20Ia7nyMaDoFqhGQFICeQHxEo49zP0mFKxiieLlA84ZKGN+4HgiarMEcEXH1g1kv66sx4
cILAuPlw+A0faHj/naanDfQTV9fV3OEgA9QWMHczILEcSSIZeNyHJaf5L10V4C4N0I4cs7btcmqN
rWchR1XY767KpLrmLLVRimYYu6b5CtNSA6iBSv8+QXg8QOAzqo+CjRil0Jpst8p0/3C9hdndiZq/
scRSczjfE8VZbPf7l4FWu4O94/oP+3TtKzY0JtwVfGt+90epWXa3CqNa959nWsg8ZtHEhmuo9CgI
pAMFZd8Hm+26a9D5PMg/n2a/fq6J5vJz/H82+0AdCKtJPa1RopbrjMFWQmflLUdTYQKi9MRhj+Qt
sh5MtLkU1Izq03wLhIuA2Rk6VNsriYjpbnxfTvmtxRWEK/sAzBr/DwSdOY7Zn7L5X2SpqKAIU/29
Y1/rKSVOqxUhbTUtVCgVaUaQtSZs5+A5hSih1Xl8PtdwKcPdHPxa82wbiUTu0TZKj//Sy1aCfBBY
BzNoEdgd9t2IU3aKmDJG4EB7WY42b3tsmj3kH3qWf0Lfg1/1+87VD1dWioLn+AT1L1vN9bqP+K29
Z28pwnjLVL77jOFGatx5AJQnmcov4lWmoPBRyUZ/lY2yKc7dA3NoM5gOsfPFao0lZT8HVfr/qClq
IaVuUQxKQpzzESqa4682eZeJDuEL4SExjPn2IcidWYXSMYb6Jyu7FNuuvSX+MEvl+mbbfO+PI+63
AYs5uup1P3c24KGgAVUOcxFJU7c7VO6bt9OoNjd75+ogvkM5O3HK+dQ9+jkzQpQoBYklDbV2vjk+
iCqP5jq+hfeOv0S+l5mZ8cj4QC4bp9CFPISZ6qbDRyy2FQc5oVDqK3FyLQOin/QPDH+vOYLMc2q8
SJyrTaVv5A2HUonojlFOnJKvnEUDTtfqTiUyLSZvSS1U6uuvHEFhhYDuztAmDS8mJb/13perYwZC
M0Fhm7twLEfp9vXpU4aZ/KhT0AXN84vI7FCF7KjTNWO3HclyyvetIO/0jBaUWUDwUu6MJqxvPinw
NomBI+on93d9lQro1mMCeN/uRoCubbzrbky/W/d3X8tXtWetux3/pAVJejnoPrpXoeWmUHQUGc8c
cak34CscdwEcuDrHR5tM3xKqpf+jfOjPI24DjhCy9Yw01pg7WKZImZ5v0PseGLyPMHHcIzEei2Ny
pPOgIujNxTghKTW10BYvU6ScHbioUwTvzydBaD19cK3T4xzga3ix+eE1xscgsC1I9fSRN/Xf2bQG
Dl3PFuiv+u3BuDzceOFoVizxzKXWoooJsGaD7cNsDDMnhJOLnXCccTTh9Cs1YqpSRc3KL8FnbX+i
W0bcxMocNDdHfzhw9jJFUD/Q/z3TZm+7uTEReoV/1ruiCfODuGQ92K4nBOjTrGHgzgb41W8Ld82V
B9vQ9oPX8685P5ncB+yMJw+OIhPfk8HLb5Xrfd4zj1WK1615HZGpXVQ1p70caZLJzvIhpca4N3P8
KDO4HeS+U0N5T58s/0XXOYguRbzrfqIP+kPMufb4ccsjq2p0iiHrOkTPVQT2Y8TIhyoPIsieWvBI
3GH0R0PlJUYxUSIb+ySbfzXPO5SyWg2L1UGZPqK/KOnqpJ3Dy9Dh3XE2K56fov6rbgbUtS9XUAHm
eUSInpauG3p7c2oZejJ4uQQ0U7T86wNCYKnpmjkzTSvYjR+xGYWREU4aAoNOiJTtikav+2iM3Vy5
1E9BNRfcc/l5di5NiDfe81HX/1o5XjXADhd9XrKSE9dLGFeV9BdOMB3f4kxUlsImh5WFSTw167jO
MlUsiOPvcy7120lbwMl1BQPM6p7SNlptzVX5+l+mfqgY5vg5PkoCJI3QcCBN1esKX28SwOJaDpWg
1qcCgNC6h7HbSLT2mxbB99QNXZ1AWISSjzlwZCLYJwfC03AOWV//2DQj38GSWQmMr1cGMRWYl4KO
cTiaNcHJlTiIdXsYHjxwsVs/Xskv/mguL1YMoT1O19mVExaQTYyk5Qcs7lma1SwcXPYcQ/7oAriO
/RZTUzQdFm233yOxBWqu4RYLhIemRPFoLSS/PKF0fR/5LSo2RB8TdSSxTbmwFDA+ZDzTOaTvcFkK
FMNH53XO63267AAm7V3GTkgdWnG9qcktvnYkzQ+BJmap5kvld+NJVsA+EmquNp07EgVFgcBe1DRd
I2+RNRi7kZMvaR6d7tPG1Wrs3T4rHirtD73z6C0vR95sA6o+ctRxIY2bzuY1TaOam4h53Hb5NfLV
qCDs9FxvVjWuBRVnbnYrxGyMlnVZl87+MpgK0ZGJffN1JGq2IeBwLKuKB3RiAHauKf9TslBi1azI
wzS4kU7JjTpwxxv9Xt7O8e4SEUkKI3/BQCVB5bDSD0ooVpJwha8pZekHUFA6uAHhqKAV8SGf7eq3
NwRZ5UT8gDJ40z2sUjO3YPYyr7ocsrt/35b3mdvH/l3aSncRqu5S9CUdBC1KFYtFtY7LyTWPLxIE
0+eRZAPF7pTC0oyqnPL8iNtsHOdcI+mS2dEVjcqcc+LH1WiGjpDV3UfdrZSoGpSjsHdmVAynb8/h
6ItZ1KMbl3CHuaQjutQZgGKMrg2GNMGdm6A0Hja7FNbCEjmZwYUKn7No6BpmKLU2VDyFc/nrdOEg
KIHd0CoytBAWVaTg67CWQLvtUJ0l9l1Of20ENR7N5k9eBz+bJL9W1dwoxruFWDip8JfNAhqPT/Jq
nFFWR9QdkWK2XZvvLPXhDIGLV6dPfWjsM4tLJyPswQb05+mp5aiCwg7vhmDlo+SY0iAHeSJeeecc
cVTDWmCBf5FyYunYysRd0IBRqNK4XttMWuLOpJdmOVIrKRazlzYm0/WkfbavsHEo4XGtl4LijLeZ
nTSnb/y1vTic/VDjhICV+zUJdJ8v/4mj9P4SQMvBWmbhe2+s5X3TuJFDtgQO4DcEuMkYAO6nEsWL
Np4XQsKO8bCfjqsyuM/QBn5VjeckHke3XIdyyWzxLYFwIEovqXYI1FO/nalD0Q0bJd9tc1yOSNXV
JluYOVwnJVW2ENY9kBPyWLl3wyFxC55rgxCKuyuIQvt//Xr0yO7DTVuD6r0zc8HCMtnlMeUiMFmU
mN/82xzfbSrao1BXXfBiinaoWeiJbZDFC94gjlo/G/PHJ2ZcqLVj4SAdd6zSEQVVPjWLVtAhhOWM
L1Io1+APukwDpZBepQtd60TAOEGXpCff+IqdbxfSsCrjVOiVLi+FriaJsRdM6i3OGx7c1g1jU1ab
9C6gD63/Xp15bQ0DXICaLB5PXk6CFGQK/sXw4PaEbNpinf/zqIrrF8fiMBlL9TcDmtowJc/31YU2
VuBQzqK0Ew2Utxno1v0j+kmRpEUt5SgIF+IAccN/k4p/bVhCNopL/x+MxpiHB4zzmeoRvSZ3xOsR
8EMaXMH59pbR3WniHjyDRVuZak+CvdCtEO+ANSCNPJtvcnV/vfMkk7A1gbChFs1etiNjoudDGL1G
ttCuTPXtkPNXXyLSY3P7GrMXxau5Mq64ZvNDFOwhp0Ndiy1qZDZqYYDk32PnmOPIRwZGZc1zOimA
llG49JDNzAYsyUN6pPqK7yXwEo1FjuBpM8LhgDVx9ZNrl7Z1K/S4+pvbFCHtaxxiHqow64hFn3VJ
mwLZF4GiYwvnnZAwKsE+74UkCM+4KgfmfSPd//KRIdTPA4OBc+MyGLWLaddHhYJlNqKq4VIeborG
sLapFM/O/wc4IelZO6PSSniIP1UEHXzhp+5JMTEQ7iwoMoeZjbc9/prkkBz5oOW4Edl5Z0oL+8a7
3eoGntzQAZBRLK4yOe/u6tvhogeNjMxCEboSgj8XU+rn/raDjJlwE+ix8YDc2AgvjbSjmvzxRqXO
w3zZcRMcerbfvAo0FXoRxxvo7iT2mHLZbc/PZndbmY441Bq0d72nFCjTI2I1RYAyaudALmvYJ8mD
ic4UV5puEQpWXEFzDGeqXk+p4XaLWbnPDjE/UlgEMn3qMKM2uqIo+P5KFE5KYU7OrSHnqCXlJZeU
tP9yC2C9eJP514px/0lOStbcgddSt2d1GfLuGiWS80CLXmtCPEEtJoL126UnmMomsILGf3xsbcAa
1IMljCC9JiokOOHf6HAdh+DttknTpWo8WkjHd6XQaWDws95gPB/owNoz3VLi/T2218U+sikvce/I
tFjKXCNScGef0GXNx5zT1QLADnTVuJk0YLIe/tH0aykgyP0BouZaWHakQ8r5u8hlKYEohiwEbVa5
6sZW2jz8KUGrDZC3y0vQ6IfbBaBgT32ErjKWSRVfohdMMrY0lkTJCc8a43iGI8UcfgkHxcedliqK
T0b8zTbtuUzmk+Lp8Sce5KNlnIkKAgTj8SeiZI0OhO48V/2Yy6Hsd7SDWqYvTXuoab0DJ2zU5SAM
lgQ2sR+RAWQUZbi+SpLkdSWb/S+cqprHW2YsDHh5w1lNjzBS/CiwWgZT2rz/gxdHVk3Nc/FAFuTP
fDg84nV0iZaHCw7wkeIzXtkCeYdzQCzANv+lZz+aHlBMTgpkyGw6Ao19LaiDRBDVecQIcABgl8E+
E+4sN25aYXGO1FuQVof/MEOH+rxq/69A4ZJ8O874cmScY9nsh1qRrlFIte27PjV9WuT59N9ZUrde
6zwIdVgVpDk/3N4dqJEYXiOQGAOSNcAvE7EPVbm+eEZDRYUxObBQBQWx0a53hLIEg3vu3PjM/iaS
NznVIyVwtuZYZEgnKAvX4FCQCLdKqMKPpWaKHWRE+kI2Le1rVLFMtIxHGOGS0Pq5w6dcgoH0FKa3
JjkyFEVaxdtWgEl4oqrMOePaau2hEU0M8gW+drVwjyJ9m7tLIxM1J+kFX8kz5obIe0Y7++vHnHmR
9Zj79n8hZJIWi1tf1ZT36THFOLdwv9Dsvmn4fLR2TKUl3/QkmExxj9rVfefEeaASbThYpryRW9zf
eXlKARsmgQ3ya1f1oHYb8QypglEqH4i+MfGRiugTdrAT/FD2Qpz1QtQjPz9zpnAsq9wtIaBQ2oy3
/ToyB86xnFAUrIPtVLW7MEgTrHoWOQOid7/6CpsImNzBh1MJ8FKaPCwwG+itZegN9a+yAnM9GNzv
366KwDLCSXEwxkocjUm5fBkG5gIk4zgbLhqN2n3MhH0jbncHPd5c5rYfOXaVrItFnHV84hANAnNl
kU8UN0ijz88tGi92nouYx2gMhaSIniVuuGKOtF2GJVP7EajO5DyU+51Z1Y9eGMVMDsd4CiLkXaBM
H3xY3jYzJtNTX71m6BoBVnB44YfzFHXDnqVKt9ZxT8+D8gfZ2srrewCgAgW2+bQWMq/RFFlGLSLT
x3IYilTySuouLD6EJsf6KtTCDTPKPMIvykpkx3e2Vye9bdVtPaxJkj4oQ3XGsY96Cm/VPk0e6Ps0
OOQSPirUdO7Rrem0Jp4gFKLhUvhIjXix1tCM6BOxQdhzFS17ioYqszWHteHR5Jgz4jM8aTyfuzbn
3IFKU2RuGmgZ6NftPdT5Ehm9Q52gsjCGtUiWf9GDvt3rnurPCOB4idnnqaC4ilLsJT5najb36jlS
IiHrpKU4Ce4zq0eJQIML/lzLCxaJg4N/3FghG69NroTCLNUsAuQOrxyo/EmEAJk5sWNF4XJGpMJR
+ec3zMDDzUT1t5b5bdS7DqsA2xLI9Me6SVhVNxTSvPjaZKZyxLCw7Vww+ntWQAES6qOXspql2LoS
BVuGpFtRSXq8bq54pc9x1hHrq0Dt9e+99Nt4tWJE9z2XBccn/DdYCePYvriKrnjpsU8UeLNV5nS7
wJGEXyOsRsZNAHQFWngcn9/JEH9BWcftSPZylNmzv9MaoDcI4d8jiP5Z1hHQ1jpaOUGQ7VDpOPmB
WZeAOwLIBZrpWTg3YyJoqlEORpx4u1Ylx0M6WTItYYp8rSA1rGep1dFqDpthQjcFjaZZWJSXMzhk
6OVENPv9bEygWMbN70I9n+ZqHszHi+GbzFMf8UBW4SDkrKYlVt4QkCEoimgupl/URuEsg5CSuMmG
C4CBmkXTlXqA+lbOV161Ab2W40e/XTANsBPDKBX3s7cutRaMOqVHwmgWPCzC5wzH63FpNMFwR07+
75BpHFhWlO3GnPDKq2j8OmaOn2ai+BpdD4gsL7gBNgmdkG9lwdWzJ1dmIUsO33XIaePKN4d+ZU6u
QbVaD26W/oYU/tJ7yi/LezJrhLu4AUEz2N7+/hRZVXq/hloc3c63U9k47WxFpgxvIYAQ5TqeIwXk
3eaG4IB7MilYxshsTjz5kRw/lyD6BzgrUwWP+WNtOcjWGcCHNP+aECrzlqict+QKo5mH38+KniVN
Falsh9GUmf9dRVA/NiHrCo1l/CGe9sq7BtT+xXjelez/yPIGzcWldZiFcwjBDx5Z4haE8P4SnpJB
i5dkjy6qHIInFdJhJvQv/RJ1YCdQVBLxRHU1dK2PtfXRNRwFhmc9A033wOz5ioToAIVnvcIjLo85
E6GQWjv1al/BdGBGBLPClM0KNcwabMkN2yDNZFgx5SmifSTlmEUdMtwEU3hdrqf+XqzsDbODqV5h
4EbvOAXsFPzLKU4cluLbmyxD6FqLezWhCL6Nby43GW1kCwGX7wik1RY8Nca11kZ5n3JZ39V4P088
1RcxHknzdFcVm5UDtN8bVmyZ12vgWY9U/XlRdwNm2Z1e+Hd8WZ+esq+ZZMCcgInwNcQz4BT3iojL
p9CqUddppeLjVLb0mA5R0cltjWDpqHRts/1MUsfnZJJVuNyLUpGty5dDsthekn7DZCwcJ1hJz3xo
dbrZcm/Jq0r/qBVMcKxQ0TaTuBpyfCNvSaIJyMbVh+gjBvAsj2crNIhfOa3lI0lLAXDhiBCWosQH
ACaWlgt9sYZt10t5y8cfuHTFCtF90NbLHqCtSQw+AuLP1jfMCk7Ya35sFAp82EIfiV1I/vByvqYp
NvLSvziJBRLbe5M56YU3YfWJQkgbPxxz7L6KlcgtiVAaPKqxWb8CWvrOqGRvZ8haahWbA7EOcbLn
uyV3dLtehEj1AHDyrfgbQMqZeiQWrIFqMkub7LsYDT3ujhbC6/dtWOlmN2qUz3rY4B3kXNrjzxFn
bAmudxkkwtRblkDOBy80FeTLJy1ncO0XD1K9buUVFDaHadLhA+EO4iO8YIN9dSsI+zz7oIDlx6aQ
xP+odcGlQA4l+PAOdjIa8Xeom2/8r5g7j1/GwUorNCMl3WVIpkYQ24AZx8rJ61jj4m4FCoNC+HTN
/jcOl9t/cu9meZl9MVs4hlpkvERlbo9BmfPI5DK3d+zoKq2Uq5ueE6Z7TXFlSpzjkPGYfQeITlgc
QzQdi2MiSvulO8WShy28rcizOeay1DtTLHkTm/O18xNcntYcwl5wQ6iUjP3x3vTFdm6+8jHwUyYH
WH7gAKQo0MVEUgUFOMBfeXhL++0zNGZgMz+vA/I6qjWKwI2IbSiiIXOtg+fAPjHqese4NArO+a7u
YfiN7zT4aEep0ZPrK3rO6KJtj3MJTe+ArncfchnVrHFjo3KZ4q9W+oSJj9v/ez8FR5Sv7a3EmiI2
TcLwjE2/vkZ3f+WPO8rpK0Apcmi40iIk+GLkMQN+I2EfmvspnBGr26Q7Uh0quvHluRynHfaQOs+r
k2Mkh46iPcfOoauseVfs2HLmQvnMbIvGtQWICTHHpyJNC2b/IvDcL8j1S5fMu4/3OZc599KsTkME
2M6dauGyB8O1ycvpXUBnGS1UwBFOdSKE9JKMbgnQDVXLoJU9TDPCMHI0A6Krjstjme+Yh5XLAhWo
j/px+Xj2sGhRXFHFCMRERz0hIXwNids8Mam/aGNTlEROE5FbBg3UR1yQyrLmGZK5gaUXFouY8W/K
jKs75d+fYzlQXSgZ9qi+7TxPDDkPJa7UeoQGRAopwW5iM2DeRea+RESD8UxJhJSqpPRQwXNiCe3v
jZ5qjlhconWx4Wql43P5sBrAJ/zMUHWVwZ+CtrVj0Yl6t04sUIOxVF5/6cIZrTLeR1eEfNkDf0HR
OkxK1wHumB+06jQFwLamO/FYpR7iCpQxlxfMPHtbqLwmtUnov0npCbgIfjpwcJDK3yaHz6XqNbKV
3d/dICufFcWgC0qOM8hIXvTe0SYihJdzakczSaRSkOtfdiBQxw+Agfo1J+9nCPRyyqHTSmEEH/j+
A1Y5Q8yoF/8U7GMDzdn7XCotJSX96fcD2liCfKgt9BFOevXd9/tYFC65ValEt+l8vP3UaBqzScar
0Skf4z2f0qpSTI//mOUx/N0oBMIf64gVpE5Ay5x7m3O4h8qNFaLSS0VoDT0B89fVg0+eWoUu4nlG
i/BIBcCJzXNWbZtFobu8gXDOQxW+Bb3lomFPvIlrBsnxQ5HjlwjBvWcNM6OY4w6cZzzCzEvtwodg
22Ugpqzou0NW8cbdo8R1sWN+SsxbaQw9UmKUf0uRe0fVyQSKqRY1rwsDM0Ft/uSRFo9Io8MRGGBj
WgRWOZgdUCopX/1DX25tnJeokQinm2ltXTnmrMtw1pqz/KHDNWqESUmreyWW23B5JwqUfRROYbXs
T/x2/l1C59LsSn4gTdsN6xRX/AxxW/Y22EslRP9zpnEFZ0ksy2cD3YlOPVpRy0ISAqC1nrXdV8y7
qNeKmU7p/rNHB0S/Z3fTjwchSgWbg8c9N7cvssnOZnQi5LKfY07se5uSpRsGJ5GqxThEmATDVmos
+xdXy9kW23ImiVMsYfC4LtVGt48oTnvBgAbAr8SUQqjHazHH8AUyW6zMPelmenjAuyk99QV66Zn1
xQbHMVsVEzPZ53+7n6J46FAJiPnMbKuNIL/NayTUax4a
`protect end_protected
