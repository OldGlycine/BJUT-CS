library verilog;
use verilog.vl_types.all;
entity npc_tb is
end npc_tb;
