library verilog;
use verilog.vl_types.all;
entity D_FF_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        QN              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end D_FF_vlg_check_tst;
