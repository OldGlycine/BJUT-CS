library verilog;
use verilog.vl_types.all;
entity counter_top_vlg_vec_tst is
end counter_top_vlg_vec_tst;
