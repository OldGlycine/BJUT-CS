library verilog;
use verilog.vl_types.all;
entity frequency_divider_vlg_vec_tst is
end frequency_divider_vlg_vec_tst;
