library verilog;
use verilog.vl_types.all;
entity expand_task_vlg_vec_tst is
end expand_task_vlg_vec_tst;
