library verilog;
use verilog.vl_types.all;
entity D_vlg_check_tst is
    port(
        LED1            : in     vl_logic;
        LED2            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end D_vlg_check_tst;
