library verilog;
use verilog.vl_types.all;
entity reg_N_vlg_vec_tst is
end reg_N_vlg_vec_tst;
