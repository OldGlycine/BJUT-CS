library verilog;
use verilog.vl_types.all;
entity gpr_tb is
end gpr_tb;
