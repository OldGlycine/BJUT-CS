library verilog;
use verilog.vl_types.all;
entity dm_tb is
end dm_tb;
