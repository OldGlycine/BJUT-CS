library verilog;
use verilog.vl_types.all;
entity ifu_testbench is
end ifu_testbench;
