library verilog;
use verilog.vl_types.all;
entity seqdet_vlg_vec_tst is
end seqdet_vlg_vec_tst;
