`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JyzzRYOPvALd1+n0h6OhFLeJWpZqai+m9G1gTt1+XdvmSl8CM8+DESDkmdo/iSod4UV7qKGdzREk
xhurZL7CdA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Uh3HQ9MYQCOnfgfbo0Xs+fYfRhBW7I6lM6nFARWXzDWJdbXLdQDXYmHQftz1C1OLUQQE7C4dUBXq
dT00dZogf4QehqG4RWPk6d7F3tn7Y75QCE0Hwxa6uqjs7+oXdQh65YYvgBS5EKqouNQgbBWirj2A
/O6p3Dk3LXi1PDC7sQ4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
b03Avj+lw247JKbbtrBPcXCg9zTXOiu8jwj1jF3NjD1nO9GHqik84DfX0V58lqrsrH0D+SmqG4qs
ZDsMe6f9LVCTEnKWmYthPlt9PzVWNYgDu6L6HesLNnRMV9TjJ/scQsgpJN8+vWZSpWvbmzJa4V5/
YDFQAUnzZN4qlNwPAYykHK+zBkPF2e9FhnRcpGZL4OYtDTLMY0EDdOYsRLxL+5sELUgEdaIZNLVt
5nK+WNStkO1LGCDby8DvvdpJtFQVJIrmH5/ZqUcp+qSSoiyx85R/9j2BwYYfh5iQMUgbKoJOVJpl
AwOZ6sQzKTlp5Jo9k7AJXzWasteEYtt1y2LrcQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dZgv5mGQWdpc0b+WNxvFkdblBIFCaMTgSCbDL6OPVir/NIFh2mbMpEDlagVKrhDqtUspl2WJUIvK
WVCPokONeoUQUX2YXU/2M6cJDMwC9P0Cta9LirDQcX+m9xLP4zUi6s6d2phb20vdT7exxgjE27i/
OiMCLmraNlYn3IoSn6WxMekR9xOwc6NwqOntFAL8EPrhs2mFUXBlDxxGUDMmRoSX3KAf1Yljpkq1
ElzH13NNaQAj8EwskvhUKS06GtHycaKS0PJI6BoqZfR8wmI6OLlnwaBnwBU1OexxsuJZqD4RpnV/
AtyK2U9g8WHHDknhaF7VrWI03dPT+QRjMi2HTg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rGXoZHxEO9Sud7P1xF0JTgZMXtKljokTOQnslaFqfRTOADB2sm5nTbILbXiltCqL1pe3cX4d94Sk
hrk5vUjtSQvqWbw7xf+zcJNMMCTjilITlhm8G03/LWTrsTqgRt8HrZdU+IC6OfIUepPii7PxiHNh
LSn3VdihGfW2lp+slugMVUgGhwaAcblMBx9ti6RsCd3s5Cb4HQk5v6vch3DiAY5nxOR9DJupzHSf
5GPg7NkhFZ4zURPoH59I7BKfTTajBiQtJpQ3hL5INjQgkXuEonEgqG1GCqWtIhgc+RMEM17xgyxT
z8LRfywYV7oG66kJ7LM7+8ZeYA7iE7OC5ZR7cQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pFWUSIOr/mjqQ/PncvQ9tWAvzGUR0DluRbBMvWIA7v2v0EJSSwnYhoaiAfEa68QQ64JJWT1n47jd
yiDijsjOmFtJUeMTIbdZh/G2f1y71CaxbIPYCemOdxRf0RG53R1jYD+fpC9nHJTFNthGKbZV5FX+
Y2OeUQ85RLl/kbY+d04=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UcEibmP3nx2gTMiM13z/i1fcD0mpE0oSpX4V73bMBV4RliRtcJpTK9bJsaH8pNKFxCIffkbWSF83
bl4CMGv63U0uDX+XJnOXqBkNH38mqh3WF9bOqwyETCVmEfkjWqeWxwnq7Of5JY7xuUwX6hqf78Sy
YjyiaBwhQcFiwyxfeheXGDNCAxLDxKUe9RJLUilmwCUXjHTTFKzPIU6/TYxmMvhlhSgZU4iWRNSu
6T3hrxHvHM3h3FEsvqNIwCzPVIVfAS7ZURK8qWlUz3TipTnEiACdWQ6rhMUN+JygWCHp36uogquR
oUhba41/v/CLPaJ9RrBJUItxOGKAjzptwAB3Zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23056)
`protect data_block
q0tU4mad+YgA3IveMt8gJXoqoM24JjkEqHVY77WGT+BacebNhl+/o3wqq1DPzgFNCjJ4zVg00O1O
NpL0eyeYuabvw/H1xuWHw3TEQnDf5rtzQfvZuXxZ98jdBwSELh6IZ4xNXLAvbnevczIBLR18CrXB
vBwVswwqvBxNpRpQRXnrzEEk72zW6cSbQFo4YnfpWVRjF2M1qGKTe+pEwKY66O0LCJ+akGOpzMLi
Lh2DHkPJUCU/Eu20yL9V280+OXKwRm033C6fT7oCGJ4+lUtIR2CazL9aMU0r2v8IZ0o2EtonP+l2
rLYUVuypnCbyjRryyJZ29GPkIPejJCX7EfB9UG1yXi6MsMACruNoviRkR1iZmejnuPSjIBll9VtD
NCVyUE4n8cTV01an8K7tLwkserYoO60OGkPmbGfqTdE2neaWeSrWJoyKpDbcy+BzijT1AIpLk3OT
EX6yte9gGdrePHF2UvrL+YpAnTcD8dCs2aXnc7Jm2ycyR8LH7iRxjB6c6bAu0zDKwOn6H4BGi/+4
+DjlPTG+EJiyd6qDNri/2XfyfvO63Pe5N1cmRxa4ZUhjL6MZkhe/rYqJQTY0Hts/K3VqKP61+XxZ
zPjCxtmKCKFiKKb/SESAmzzP9ksKCuEAndFa0EIx0rSpwCq7nK85+ykBAwS6v9FCiZ/eC3Erts5o
/jjvZgg6Qdaygw+CYfngAhe91+sqA3Ncspdk/TMmnhlHkx0tzN5odByViFZncP7PRfuxAw3CF9LP
Gmy/pCVkvaxCwwK9sl6ILZaecqa3cGdwqul/Addz1YrwoG6dq13jbX6wYpd9aPikDHH0MlyZ5Jc+
BSkj1fx3glmErhx4FYGEZzuL7P7KdKoYaIbYYPeuG6M275BffEZE2VijxjRBVyjP3vfvpEq/Gi2X
YaDOz4vMHB/GXwWfWZfWpdu2v2UAk6W6llysAXLddDIhHO80vL/zGBfNp00grhOfogdS1Q0S6jor
PGSgpf0M1PIglvk3H32JD9Spm7Gn8JL9f7iInrhHRMEVZ3KoFtf3p5JKmnHyhbcdSLFurqvjlUC0
aBmIiP6aUCeUmxwJ/lwLUSDBf9C7VqZqxdp6rWBD+Q7jajtL384WNfGtm2/I/S+HK9n6u0B46RH5
MLPwAVe2CBAiHUDl8uUYmaaVHZrk0VZT9Z08i1mSJOGJpU6zSSh571O/Etd8lWtcw3+o89M1oDrb
+DfA6TAdSj2KGOdvnD29kpVODmTYywaBlqs0KUmAnl3LfGt3J44/4RzNdlXo96e0f5fl3iWA+ZD8
RdySYSsN2kNKe+mewxtmbLVQpKxvJLBbwEZu5+EK9+klK5bEeHL0UkSavvrxC35YzLKOjcUQQjj0
VAVs/1z4QgYxyIp0RKXYJxwkp8PbMWX/3KqvkCqVgJTNu9IAm0Milsixf25tCqD2ssgSSN/yS7D1
pzRwOrG3j7yn2yVSFMQBrc0DiRNRLi7p/kUAw3blKT7NfvJiO/reQQzJYsgkVv4wLyfH+BE8dTMy
RckmLejZiYNQkqL8+84g5bckQRRyp0Qf3gzXJ5Woro3CqUxQ0EadWCUaKE1UFYDLwnATirxFPW5/
PzHM3PZCuv2tH6+PtXyoO9TEhl85fhUi6lGexbFz6gPtjfpWcVZ/1P8vO+1H8BUhzkXI+D/zhx1y
hrE8THdfjdz2SEGsk3x72uToppOhgHNcmHlq3hsP4yiIXaYWGIqqEK7mYTuIZxkocEWQCJW5wtw5
LjRMaEfKLP9c8mOeP9V8eygU4PDtigARW3sUijsub7co0SBQPOBeXmQK7TZx7CDMPK4g26ulTOkg
0RbkCsmUSvEXldejYfFbDwwwwwlM4nbMWDz/wYfJc4S6/DTNJoCFT3VD48abNBDIyyrMbY6harHk
F3XhlGC5lAIl2hdFE3tW9Wz4++Z77ew6RwLqZY5WG1ywbSh8LiPrkc8m8GcQ4+eUo0on+gkKzu7a
K/fTPnos4/L5LDVHNCLK1he9Qa01Rr2Wxj1Cr/wU00ShfvbMPO84ly/nQb+dZD9zbW2mch/g7LVP
g2m9gfVrN/7kuclZMXgpTs7U8CZEoHdIC0m1Rpz2e7k+vMNf63ExwGSyd7997/rdbUKYdymnEbPC
he0XKuWepv0614OIWAMyVB8oFH3Li06q0v+zwYybGcSkeRwCr6s5OP5VS22qzIgt/8lYMNI1hDiQ
xIO7LUuZwDj2j2pAw4GPR0geqiA3QL+AoIBP5fexfxbuVjnL4qJaKxFIy9ZEVNn+TA7X9eW/1uRO
WB9PyV5Gq3i3am3qfZ55AtTvV9Ja1gKjV+l/CpO9sxFoxNGMYyVSAzKDGODU1WUbn/tHezCcykx0
JQg4Fm9EOpZQTok0tn4Eo4Ks/W6YeksUfB0ABBUDL7Q1RgrO6zhcMTt+/Eu358dG+zmFVoSexJMQ
J0h2M74UP8b4OF/yOewmXe2c6nXL6AhHEPTuWkMqNl1f4q0r7uCqkbnezoCEPTxyviRTHaew648V
QKWLd+Y53yyXVFvtXhap29RzYTVRZkGCRlyZaErs+/A0PDa3xnu4BX3TBzm+8HU7CjRY1HnGlasd
daYnLZpdAyHyaeCw5awD7jnNXRLSqL/4eEMHN/ffZ/5PvdlH6SjpORBu4j99zvxeP84IaWWyFo1Z
KiD0+t0K9Ezp+u5DkIRHSNe1idl+6ElsaKQ9qZTY1ML36V8QHfsbGY7UzHAdIdGuPHGhhRU4bHPy
ZdEHtqPiJAYfEm/EUidrUlurdXlTYGk26R3423uGJV/+J5CaUVAdaFeZcwn/sjtehiqSRJDIR+fN
4bQUSZknC0l2NDzBW8Do+s+mgttCDg4qhQsXUJQ+yzdeXG4sBHVVLjoYtVXXg9fKbOvtwa58ltr2
YSSaU6C0/Bdh0Tm9IQCct4HxNBo40sK8sJqwGubMI/Dx+A6zqdijlyDMAMqcN9xj3mm4nHBWbDYW
kO6bDgt+5HjNoVLPXHBvWafaaAK+9Kckrso3Nv/LdXdCXCksh9l9XX2hp6SvTCia40Eg16Gxvoyg
nKvLfm4SsnhSJ0RbPbecyDRE9lHK0kZ0jgxanDCdPT5sN8LkFuQiejpm+yLQuoFJtrU8CIJzGKMo
JaIQTIwmFg0pQnKhsqhlkPTNn0m8+r6ZRJVsPecxqXu/hJNxNmTP/gG0g+RVdg+89AZUDj6lejyU
AohwTBjas1ob9UaVJm3USie4XJ9/vl8RRO6RCny+3X4xp1qvOOzDzMO4BfiVxhW+HQ0x67Oo4yUA
X6PrfrbC6Oqa9Zh2jJqO/AGLKOK04vpitR6Y7VvcbYWh/TsXF0os4lk3SpfPQmaLkTbNcAJOqT2x
6T/cqmMb3ljXyniNaMfYDsoKvjZgK+j8zJibLSoEx88c96Iar849mo8NT5dzY69vZRvG4ObjYoPj
vXLZmVJXWDssRqEyCOJmRms3EiSOLUduh/cDnq05s9Vz+Ri91NkiUUK9GxSzLBW3CB92pHLXL3YH
/kjGOa3eTRiyNqVKn1cxsGDolp+fIt5I+gJZ7/ftqkn4Z4S71Seu3X/TJrOqZWzURQ3q7eyUURWR
YPKHdjUCERknv6Mb/p+4ozFADdzXZGOFhlbWO1A8ewixJrzR9Bkliq2+c+ztm3Ymmx2PXDQ+ZuSu
xfMuG5u5ySR1bNSJmqa3z1xul8PzxxcpPOpZYOQUA+swDIZL0PUVNihKwiKpOPxZn/off2xUw8zS
LJUC+Q6n7qIGykeBKW0fYYDEDBi6brBbWkZFALKblg9EIUblNU0D/wtlxo058mWQl1gcqWMqPfQc
/j7034qG/zg7MfDJsAqBCfiKJBI3CjfORiSJKqmWW5kTRmmWS8vNjfxPwo+jI398ltuPjXINK2C+
8HThZidpvT6v+p4/uqHPYF0DQVrDVELdW3a5cpnwHs406eBY/EDnXPZG+4WrqKZve2/FR9HFFZvt
/rP+wMmftFUIp1y3G74CYXum/gjYAXxxrfiRZmuaQO1ENPDdMxJsKQwRj/gxqyu/1ZJDLBSFAhlZ
0Hb5tBymQSFkVlplBT08osi0YuJHlNKD390k9EvXKKhtC1arRP+ybltnWU/b9MAV31PqNEIYE9if
Vi8F1VzeMYqF5/A59NzC6H3ZNOb/JoDo9Yw8vfPTOLrYo34uU8xwLntgMhto9gXREuwDq/UkuMQc
hgHvi3ld3b7nGlzo/MRiQU1xQBE5zj8lqIMf1x81Awlj5yjH/pq8VOJg2UG/nCSeDaBeCoarzznD
grS8nljBW0ug4RzciHJSg+/yxCiF3JXsX4xYohOo7G8nQ4MDaB0LRnES4O6L0mZ06aRLEszT5vDX
jN8hMwfykOvlthadsnBNgqvpr4cTgFLlvUyWh0HFK/QBc4bWuSDFYx2WHmf7LcU9qlV1GLsfpsPb
mGQv7ClFlAhEYliQNS8dEIpD/p0JlV5WQgbk+2XI2Gm/MbxMzQz4yiyNOnxxQXj93XBxlrfJ0qK6
Uq0V8sON8XnPlMMCndkY5naMp30eACITy6iRtcCx3/mVf9jA2XCVlEiYf2bvAIKnAN1CUMmYqtGi
wmNcxnsei4sSDwfV7dkl4GDbqgBcY+Rxn6XK0clCPfFwkNdxx0lLYa2ywXg1uE535DiK6WDcNcDP
xB/+I2m89RO56hghJ1MKmqaI2iu4Mxt0VWM5MonytYPKqS2mJeYP5GP1weX8o8MxsokfdBCiAmmj
Qb224K/RIQTaD07heQS9T3eHxAg2EJiruG1dP3XRdDgVFfL3/qWPtkypG7G0fyR8IDb4wJyTI4sU
2hw0wz4aqDFoQxCah1gfMThgXKmLOBe3aS208hkJ2MKXNV9khF1nUs5U1NnC4j2p9Z+bWP9AoV7H
z4EInvR6S0B9qgZkOzDWuHOZM4JYvKu5YzTtpLqBr1A7FciMLFZ/P82qP8e57P0c3KYXvNZlvvFD
Auj8BN/iafxzK/si/UpiIQQkBOAzNtMBee/Tc7La2ruRWDV7o0J4xb6iYB2IjYuOXRXytFIpAbc6
s+k2cbacjh97F3XlCjJ7cKZpZvj2aEGTISTS/rCZCHGBFJFOqbXxu3gK6AHZTubYi02lh2v+ssTD
DoMSe8al9dlmFEDEnay9O8OQ90088koLgptMt2/WZq3YSxFnCtf3BGFt7Wawr1xh4YRhpJjByfpd
v9GMNH4e66K4N989LfNlPCYKPWUrPJV9qRHAc/BedhljUNoqwCszwulvQb+bLY0IZp5eYbqva4ZO
j+PZfqte1AH+Ymw8x99wcWLyIhEAuHWfuBkDO1KYDVTtJ1zzrPl2O8Po229rZoRQt9fXOYTKkq+6
CnsmOi0M/v1AdWMOs4qTOuT0jJSALMHieART+HaSLidybiZ5MQbcl0XhZzhFyeWGQo5sGQoMvwO5
gHdOJOgMigeImTi7sSy9usrQSkfbKlGWpz22LQR5jlJ7CHMIdvZpWx1PHUByEsfQlq1I3bCFfKTQ
ecY2UJS5rPpt2rcx/QPHTz/xIj+Viv9yIrxzEWFvDpbE5zT+h8V/PiYbZ+ZsxS0mnSXTX5US+I6z
K8tJBguVMeBm0a983h5xmLD03g44a8lnfVbR/gIC31OlA21vDKFU/xQBB58pH4chEHaoj5d4ZUix
m/hfo2nspmfXrirRV7jaql9sTJXdo2UwGaP000QJg/0cjG2gcvv3yrS356WAn1QNGj57chdkn041
TFCtygFZtpFSjWZpOtUnXQyafVbPlZ7GF68y+NU+mSDj8sKuZLTHN7d8MXdBiQkJ5lUNK5C4xzVJ
xdqNg4azuzRN5wp9WtiLByjFIFi/2dVCQ0974qfKDhpl0r3paPFSQ03moHcs4kXrNkPzxwgyFJxp
AHrkFIGKdHh1i08ef+ud9RfCTzebDz0BeZaLtOxNQjQQNNCNrEObguX5joJYUFoRnkeqtUNr5Dso
DdPzN4fSdwQKqWyyYq/h9IRUWt4XmkmNUNG4+NF1tTr7PATXZqx5Gg4pzflSmgWV/oFNxLznREUS
8dpkIoc8DGKgGtyRdh7XJG+Tzjgj1KCiSMTi95kr/AupQiCdI8o9COW963vQye+tBUHSGpzv50UP
VuXSEn7eGT+cT6WjPqKe6AFhq32H0Ec2rIV2qeZ35oNLhAAA5v+s+YIPmVGiGSTw3fzVm6so2Bjl
BKKRxYqkH/UNhlvCRzPi3UJYz3nO4nvlhCQ3ZmuE239SEUi0gAbACvl8cUpjzMuKrJknPfXIjIyr
1utJYFWXoZ5O7ACGeOD8lfqbSVfnrvnzYgmyw00U0pQ6BFcvOCjEXaiDYeBI7Vl/kDwx2QfZ6OMq
7HtixU3ImyC9kFp5I4IaKH9KC7o21ftDCraVYKXBnhhv04eijXioZfeH68F/A93QsE6kPWcoPYzo
H6Ub+hEOEaii75wx2VkiFD1TFEm94kvO9tI0dS+ng5+q1aDmF8cZhs5HFpdmpDYgyZAHBptMhJ6t
08edHDaJAsYST38bIvXNjCncZmhMuuWXcrA1dRJewQqRPqXOMuvCH/IcRvjLemmHuIaUSiiZqlg/
jbMvDI6xvzr+yvIheC55hA+gxIRR8HevPNN1gH5vqyFEw1i5a1OmywK8nVVI2kl61puFL6LXvlP+
b/QaLbtf8PHat1HfqU6gvSL6q23hGqkuzF7tMyc2GruN+OCZbswJcI8BF4gBvbXOl3Zg2dlBLSca
cql0YqrCmmiBmkFCl4VsJ6VpsHtYyayyGWYvDgU5KUYqZfEMqkuXzOBdUExk0268wn+q6FYzYDhc
4FEcQdTkKwnHetjabZp2AOSWAm4FKXXljrH5I/Lmyx9Srd93u4a8rx4xxR/hPRYxxGrBnY0tRNEY
T9/7E8UNNeFYEJbOjUyiJxkbBapzdGlKNLP8gaEef7Xmej5jyiF+4/aLOQt/xVfpWIXDwmi9cjxJ
Davk1cbmb7XsGYy9UE/PXBdUuxMKlR1j1uEwbT+pObFl/FE8RzZEX+AbuGzSir/cAo6qdeia4Q30
K6ArM9dMdsDusPYkaRpOkSAMNHbWEMY9reotaxZhx9zeujZ1SykSsQ8Xmehnz/bdWo3d7CBI9E4F
VIcezvJXyrCNFUBB32djVUuXUZ96ti616htakYKeMHBAEdtjWNIHkChwXgrVLu2L6Zb1mjNF2VY/
dapWwGIEA39ap+KW+HkIxuKnb952nUUD9auZE83iY6sNIP+LHdTMflRPJt8Szp9LJcyuAP5M4O7T
bYLr/0Um8xxnB1htHEUlcBc6YUAt4gMzgzMJqBFOp4p8MnEhEKx+Ya2xZVvv5fUMYHwFPye0lzQF
h+hK8gwapZqEPgfunqsbNCaqAD/QpYpHtVWnXu5858KDVf7MHbOloJaZCfA8eAYBuRcyN4E0ntNq
E+KM12AqxvVxlmDTRUzDMFoYCzK/zIPz4jvsVqtW1ahpZXLrNYClv++gjzD14LODexvz86kDEifT
SqqIDgGylK/TAOFap5DOxiqUWHMmFVVZOlqZ7K4kFLN2kbcXiaZMozY0CbcSV7uV15RdV/tgWmSg
NNKyjWvlTFDBTk+XPwSLnN4p29oyLbWPCGveYf9tdEts+1j6IC3sqmIvJNziEhK+C92YB6UV4bsA
NfNKLw3VqaJezJeUSd5kPg+IwAX/QLTmbgAtpuBDoi5lqCrTiAQUHj2bwB8r0Sg7AMyZkctgEMre
Moye+IYpD2TPJMhpBkVsfGbyVRaKmp3bSD6fPgXdR9Ke+H2zYNjVTCSOWtNvqbH0aiRlj/o5QX7A
Xl6MVgw+03xoLhGrx/YKfzKECcIywXjoBo36GmzqvpOSVSFN9W5vuy9SotXYNZmSYjiZQZB0yC69
wBMsRfKNwTHQuItZ/TkwhLIVcrgOiXG++jvxIJFI0xRasUVN0rXfdNW+XIPYCgiKI0qRTNXFw4rE
zmt7sJRDUDvJRoGeqDJNJt7nfhJaJD5p0nEaHgvxk8QMo8Sfmd8AiXCBwuhGBwk2aNMXS4YjVxYN
sGpKMUFdZ51DT4+9P+y/Z8PROn7+badLW8ItcMYQna1SZsS6dxJtnc1eqswI8e33Wdo+rcDUJCpG
6sOiyPL/UoygvkZiITL355afXOczAx8B5z07Lespgevd+zc162UtyRC6YSvWqsy9BGLIc1/Tc4zF
kE3nmjC8zk0oqd2k4e8HLb6d/afNMX7zEcTKiW+B20l6pkajlVrL8dMi3VqI6MYTHPg90EYc01yq
GZGPUxg2IXIn+LvVtmpwCoE22ZU8U6jr2DXnjJh64dAWuTDXRynQfs7YmasDQLaIl6Dw3cumLewj
9/StJ9GUciDDfpRFfrre9SDRuQltxteuf9QPTbysb29AvoEK5/Ofh840Se7ueo9yO2JHNET5rUwO
kukNR/PDqsTICitNbHyji3GZGmMO7lIZxgxizNZFt7CEWrfIGi5hZVZJh2oFhP4+gn7jr73fe0G3
lX3c0n5sCRE/8SZBe9YZFKB/+f1FB6t/0zXpB9XaGXnfSitkeisvsIgVAUL+hCT0tCli2x778z3n
yIwlTE+sjAe+x7ZiSmmg25bRzrOGs6a51AS7jRfCj0IzPZOfb9GdjKdWfDOe7uEwwCsULzLu9EGo
J1UZ4K+OSuGuPnedyCkepjaM9UVqciC9XnAinVlrRO/tSlcP9hUoURVkDhJFx/SZhgAy9zs15KN1
KiKdO8jj41PV8pLDgkAMypY18nFdGzpYSKWYcUHoTCPSbe7olJ02SD4wC4qY6MS+UviLEvz9Ip13
CNOLU814Zd3rroBEN5a5BC6T0isA3WdbhS1AbJqGjGABslZBV62nh5SXHHZQRm1HmOyMScnnKiGL
tXedMPL33YEhw9WHRNJV+qFQJxSfdzVACe0JKRzE+bpwCozKhxhBwnqYfHw4w5HuvD9/vZeXHf56
Ud2f7X3XdAr+R4bC1+COb3lu1HAqY0EOk53VIUKQh+PKZbfM6SWJDVYkeDTJJBXRDLL5dYIKPDd7
l9fkPAayhrB/NB6BXpNhr+nZdAy04qo3dU371uTwlXXfFM4bBOzoOyNcGqdT/RXdgy27YVMEJM/x
QAhfOxOjLyxU5UFetWoA5uV/7dwvJprzOOQg8IgEZnTHjvREEMtLrJ911UtzONlcP5y4W3kNdLB6
RjNo/JT1Pbw2I6+Y5B+lvQho7/q5sBt026F58ENyeq++r3UqIaYmmD56uCMtg26EeeYWAfjiO5jZ
hnZHIjmXwusF/xcDAGLKOek+otkS1FNjo+JbJSX4NLQCXgcgmgJaoCiT2+WMpXLWnzxcGXONEnk6
wvJAol1OoqGdUzoVemxkk/D9aUNdyLRj2vpO/eTdPy2VARkM+9OjKMtOtsRo8g/8PcyZpde8HSnr
JQVXgmUMztM6n6dD+ofhEbV/ApGHAwRdnQokSXECgmWSVf26LbCnX8ipMnkrLONRYIRk0A4ZLga+
eFgi0e74rANBjmd9kCCfZmXximizmy2tpE3p+QmOH8a/ynidMw2BBfAck6cus6I1YD5/zowaNizd
EPnXOTWuFFuLNfb7jm4AWfoBr4lWfUF9vURsLvvmDwMChLjC1srnfwH4w3TE9SapLuHWP0m08pKX
id6lCfzzKvoZpElBaQhs13OhwWB1h57FAbOxUKXaYhYKTKug3tVb+YTL9hBW4oXpj0xF0Sv5tJmO
+tl9ygGI90kpfQu/CDV0vWS+R8v2Z3xXRvQFfLOiU2NdTz4ebuD8WKrhlqqJKxqftf4XtIgXef34
uZHiXnXeCsXdJjkjPfT0Z9unW7VQvmEu/FT9pg8Gll4D40evicLsJwLai9ig1knROv09/CyMdSrr
4rBTCDsaYH2UNtNSYdz4Zh2zCdB93hqQrIKyH+Q17VuyD8zquptYyqxUO3mL4hmrm+/NJVhN/WUJ
oemzgGDYBghaIfWyeVcyRTv2wFX+T+kADQTJcF0ibbYN64KDIaY2U0746zsWg3YcSi43hQed87AG
4RXdwY2F74GqB3qwhkI2xwfoVCzKzLpK3Cs6+UnsWhLKf7WvBtfuH1RO6faUXy0pqhwv+5bIrouN
i8YAPHFN6XX+u0RefyG9K53rNcMZx2V/iELxtW7X9iypbejKDNfQ9IUJ+q1Y6M3QFjYNXCripGre
xuxHdYSTVpRRGFSLacRTlXR+vbEEyhKasFmIBjzTZGY8sh+eNdwMURiioBLhEhfh2KOJeREjG64E
zhCMdbeBndhKhDOgRUX49LEtxaiCICBos4NMZTlBCt9XPGx6fTvh+uIFAbHkDZmedNohGLSAP1Oe
SA7U1rUn5CsJYhiPT8S4snFe5qPh5WPpNHo5mbRLqeYlkTsQx3c/MHQ8kiCKQ1PxhqJD9N9JWgax
xDN1j3uxQJn4rFlivgw3ytt8u/lRim9uAAziuQ3ZzbxNBj6SDD1kGZX75sUgk/lH64Mr4oEaD5Ll
IIW5c6bXGqXTLDIBx8van5ABnhwcWJDI+m2bVKJZv9Dm5/8mUcrY2f2TC/N4ZYY9fqrInGmHzyyx
DfJR6BTDfgb50Scx707cU1L34UVylgW9YBVIqzAuKnJ9YM7AtkmafD8fuov1vGh1VW+ATcgSgv9P
u0RLMQPZYES0idh1yryJRB3s4pzXQ+Ty2SGa0GFzaKRCgK//jTjmlfGggizDTErXmSOnKL8uJLSG
lWF6NNyDzPXme2vxXn73t7yN5tOhaG6m4wYmMrR+L+vi+t0MarLxdEj1lxYZg5UnLWejJPyoZvvP
vljmj7y1bp3fdRQO7DAAo4KibaETlkAVZ+xwMEns/0wFKZDOjDQhoX3E4JcVDG7LeDcql11bKqMC
WZbAeMPcPvl0p6G79FAXDEH5XJGaMu47OWVTSow31eiW22f95CLz8m0JiJQRWPHTUUcVsrJbrwbp
sPNVfx5hk2BIqgsY1Li5u4o85dOFTCmDrPKjJ2SHy3rYSBg9AY2BMfPvA36JWmyCRrKbsRf73RfN
cn8W03akQVSofkcbvLThy2hI1lluXMskqbJM3TTyklOSl3PM3JWrQT9coB6S1i+AQdlBdmxZj+L/
bslZtctzVDYHQfuWcZJVCYna+7q8DtQWb3Ll1YAFIl0z6gcrdoIQjfuoj3A5KcLFW4f6WKOTjkSM
8/HhNsvAE/JnyLiBKTrLKEJWEGJfn/sxgyKbw/Qg7ZdVjt04bYzDX7jFl58/P+a3f/6gjII9e+p1
a8NkrBXhvNDt7PuJ0N4LX9uT7WHzk8fOxCBTQDKAiNwDAzVuBQRSzG+45ZLfRUtNjLRhiLl8M1LN
Nt88NrNlPveTxCQ08ZMU6xcKg/DzgynYI++89yyoortCmM2GXs+Y0xxzS8/jBMiHr9ko31Oj3stb
hRbuEHOJgVNyvBBgA34+e2xGnMyDFkph1UnDzMTD9QNKHZPLU68WVzi0eL2w6citMQWmh1G1R9zS
nlBWgCvQNhz2jDdWHQokpT1ZtOuUzo+xOZlhU1gpavyY5YBbT3OQRQ9GQqlcNog0Zqn/ksjGrWCO
tkZ5NI54QFPcUs/vykC+byTb/bXIDagMWMDmXdgysLX1ynbF2D3UbNQRx9vV8KNxY3uh0oEYGTXc
5jb2kk2aOMHx4Oj/WVC5w7KtwDsd9T1gf1mwBrna1Py1YWHVMQk3CmjSnMtZvAceXTHcDF0ev4oW
O58tFU8YvCnVHLOd+AwVSEfmTC0fxOB4jT/eaSpKHo0rZTxZUfQxUpImslR7TguhKPfnY35Sz3BV
x1ghuLMcBk0FxeBvGbVTvGAjYC2TkeciAB2RgJtgG6Lhp9RGxb4jWdphGDkNb5MJHliCNdqTMtLU
Kxn6iU7LK5UqwMExKaW872zF7OcvMFE7qXDKtbemAaychXWO3QR+udozPLO0XMuYRjVWJ8GCm1jk
OemSDInXKQCycJhdxjG9TK77dU2Jl5ney+9/g4LUYM1cUaKT3ohGsljXKTFhunBSMoFBzvxXuZPP
DBvNUh6cHp8xhxLvTpoQBISMmqBMC7mRl1hDa3NdbyXXhU138ngFav6EDV1nFrhfClLS4ywY7TG5
H3wC+Jzas86qTxFrqXm42gQEt/hAteL7Pjtsg2I5Z3f6V/TlmtnMa+yR+s63BHkM4rXNCQG3bMom
zwJ+pnGZf8RkfBBAGZb78dhfxXq6iJcccp79bM0PR9gGMlcedGCdQzDLc0ZlHwwS1yfhszUYXvRC
Ex+0CyPyUoON5cBNcwL31XWYhJiA7hCFluf9cG+PCI5blx4F31zHAR7yVGxVtAU9J5Ann1k1wsuN
LspyUAUoLBKL1DP9SegaMgInB60NI0dDC2ZHq8lp2EHkNvnN5Ex+YPZVv6nsPd+uld1HL/D0hPYL
kIndW3uKAz+How78PbNFLtZweWdjJoQxeGwUS1uMcZWGqWsfJHX0zVNOr9/rzv30c2H4V/F/sbUO
oFq94h98NuCp+eKxfPmve4TfBiRwbQ2bnVPZHkJ+2WEPMWCApRmm65Xpomi5DD8fGB5CCkPGZPVP
sqxfw8MKCcfhooKKwZgp/QC2PRxZ8tb1tZq0HRACuyeJv81DJWWwqAP20jx6V9VYIcWOGjS+Wogi
DE3wgn94PT7UNM0GNcz8wQ1HaPrXJe4jU/wkKDvHqpkJriNOOHORPvelJAx5orAZ3aAAflgy2ImV
dTwhweQvnyql7X19xs4uG//eZuyLUTfcdzC6b7p7a129E0/Fkvag3fTwGq9cLLMG4siLZsOypO3B
iupbsYUedACsGG348HlRD1nXRTneMlmwMIjAwYYNZaL1Mo5OSVxuTyNiGkNK3DPXRTNbdKb6lUEN
S8T2mCG+5fQ4hNZf8W1+T7/dG7C3mOiad9RtT7wHJOjnQYmeh8FUm5eZcZchs6rOnEZ3XhDP9oZ2
jjWTumLPzbhrUuGgUQ8Qe2E9P9H6Sw9GNLJM5dNTlXZuyjAtGofdWc9PQPUPEQN/ZtCoaY7pM/TD
xLxTuoct5MtDH4QtJFlBGnx6H8v5CT73wPGagz0cTrqCrZW/JzGkmAv6E9IuK/Lk6hDgUPJ8xhRv
NYmOuAABTJQiyxFO550+ptT5HN3fWKGTrqTpaHYSovUzTrjB5PkjKqHpm9H92DCyQRFi6RQ1CRAZ
2xhF1iB3DxFnYI0pgRq6A3E7nr7SYLCzEnUztpkAivnQL4dq7RHiRj1dhRfJwtX0FahXJE2UKlQN
Na+xS45Wz5yljCg+MyHTWtDeTWMEsKIVmDfsHDIyhf1VAZ+KwSTFVvBTN5co9EES+PJCwKG56E4A
cdDSiBhx2hu+wk5koeVtjK3BkK2raLp7XRrq5yk9qCcXlJ73jOo2wuqsVhzQu0LwvANzo0v3JzCC
je0V8M8SKPiYnhtgyiEFupoc2hBjBd0mI6K04PLu6C2eXCXEHHuhbHcb1NjmsBoS27eXLMxsd3kW
vRnCDPez0FTmPUVIRWGPBOMkYIudPrs0TI5DkIpmJzQpZ5I2sHUE8MS3PbMrzzd5dSrpWKyrTs1G
H0XoGtZsdkgolBWXnVdYpaxWTqP6BT5bHGugXt9/Se0dWfqr9u7TXUAkYO1nwOhiSGPoVLskhFRe
FVM+DPyhsk5YhnOOsILaK8tcir8eA+ykQwjHS1o7e8WVTd8nCoJ2GPwws7VmqyRf9Jl8RZREWj8X
PY9/bp9Z7XBIKKO2SsCc1CmUTuODotFfhqeoveNgE2Wwxuxxai6QgJXTVbRsx8nlCSSdoVZP9R2O
6DMOwT0yyUCx9EG7qYWu9OmdWrthmqlFXF8Jn9Lo3H41K/KsDyDKzLJktO6OhXswnnIpcjd5dkwj
8F24boFhQb3rpiKvQnBg3/IHXEzr4DRy+bueF3pHyEeAJSVkU3OBOGpVNRo1L9LsZMk0yhqhrLv2
aMzTtppbwKnOAidN0DnE1DTG6Ijr6FwWWJg9vo5iZvAp6dzUGoKIT2noS6Wukg9I9/ppXDMwQHQ7
RjdJv78vL9b+T9k4PA7NhyGpUvH8C5OMfGPwBoMxIvEpgqUysmq10YmMll5EgTMXpBZ1fEoCdZXU
Khuxac/7OZMX1cR8ErDQGS3J1xJHja5n7IWDo8m5YBCU/URyJBNe0VE/WPGxaMykfE9/jC8bfhD6
EbdU9MzpWVyzTT0L09IUyFqtXgwkQFZoo3pYhiLbOLwek4UgInWdiUARDqMIFO7Bm8OkkZmfK6ir
IJ8dDTOLh6kyz4de9AhvFTLeXixw3YYyr2+wX0kDy5Z6k08CTBlNoe2xAopaWZfquy5v7HNTKmvO
hT0Ve0jCYEleysIu8LyylNzwprx2pK9sEPe+++TcK890B420fnRuRWCy5UTMZyyWuVfKti/LGBtS
l3Or4okMZsmE6kjsxm0Et4gYM9PDePHfUOIJUvvmPegMal6HMvvUfGwJ0gaaFZcOXpdmw62hEZZ0
xmQEnPowEC3RLHY1NTyVFalNMPuiparYsHHclEyEnd6oocoVVKc+vEJPZ/jChXJsBxa4yodzaNKF
wGlJ4jwaZ3exKi10kSlEQhgCbWqYuPh41OHO3vqnP4PhbEravQCWz1KE6NVsAqEwaRHJX2vw2m/V
X8HNOiiRFZmm/xIAMqjsyLtpRY5zdxfNZXbrMpbzqDB2dRc3N0uJ0HuxLGHvou+T6FYbnPFN5y6l
bj3fKDKy5nRboo5pVB+OvQ/K4V/Sx7CMWC0EENdYhCjLrSCLF1oiBU+pKyPMVLlLw3koxMnJuawv
dBTl9G1KW+yoIOVcO7N9eH6dqNYeFjOwpzGQmBzTBfY/QUqwrdqsiV4KutRGIJUhx/MWhf0BhmPK
OeywReoilttjkINFwzXCwhmRFAYPCfjTl4AaRsKbF6d/7sX98N5stN9weZ6BuoAqEABXtKSB97WK
xkl/51VEFPQEHuDwWphmaOxInm9u8kvOz09RTBp5kYhpc16xJ/hc0xcC6CorhH1HLCwIMAsz4ri0
FDE68cfxNdGombpjNSrK1wE31BwaZ6pJyXUZReCgHaXq8UisXrps/6qbJCfN/VGnv/llghY8FPEu
69ITtJADx6XkJbrm6s52bWg8se4t2IfvJ2IqgbYftyc9mVT5FMEpJNGLQch0BSL8CIBvPHQC2vT/
vZw3G0BNA9ErPR8dKzQnf3Zae0nYNXIe4hILBYxszFQHsrdlTpYGJTmWWz/RAPZgt89gV5UtYZ4n
LNvVYVm5U+E5RsL2IucewEFVxU24l8oHbdjc2LzOmhzQ5XSckUPbiZ/stuO7TtJacCxJKLJTO/eN
HFXw7zH7Evxpl6SDFQVoygvUGDr97h4gUkX2AbzQ+/yoZt2YrVlUf5lSlkkSDx3bk46iX9zmtzy/
ax4Qv/7FvhDRgkHmiKgDZ9/CKARQW0Ioye1tRj1DHT2AgPSjPrI6Un6yyh9S1uOkYLkA/XZMJ8FF
G5hjYK0BmkcYDjzw7bjcmidFYLN+/7Ukj0AGsJQFqTjACSeJcPeFV+UAD+lczbBd0a0KTcVnDw0y
LaT/L++V6V3upzoHedTDOmsUWC6CofM8LYDHGBimvQ+K6Il/Hw9bPDHS6ZgxvW31q+lf2e1VhmtF
lIhbjqpqTFeirgw5yEx5HZB2yabvURGROkruLjERlxCToBEfiWPulOcWf+l95/eBMS4JekavECDx
nyQV1Fm2A44TnCZQ9eVvzlKmoqaJ6UfBHPFp5nXAfNqU12LMOtnbTzSuJrXGxHCCd3Y+4egbCBsi
Vvp/R7KpC+AWn9lh8Dx/H8HEDCFqFBHM8llS0HgTaQeMz1T652qau0RMK8sl9XHrhb0iUrRHVfn+
1l3MYTW0pCU7hnrIOMwMjYg2B7mstix/OH+YTNPN5ip49oeTHUx8wLzgzL1FdC2P/Y5BtIrA2gLk
NMyKMiz4F8a1b8wJcavyK7DvIY5SgDsA6SXRMVtkzFrvz7pZfmYsv30FjJAJrzB9lX1l2Id0No5L
/iRYVtl55jeIb9D+DOzIleIYMqMvg1kF6j6Ri0u3uHpbyzVFEG5SXZIIaSYWb84kZhwIzjQ67Wsg
5c6FkcX2sS/yoh1h8UqN8K1i9ZT5rIKKlEp6CZk+X6eTz6Tsplc2ofUnw+u02RO2CjCWZMEWlYMg
GhUsHg9RSPY6HxfDDhFaogJ4+hdt6aLbkd2q468J//z6PG4P0mDxsxP16368wnMrWjFaiozdOCHi
rxsEnL7ZVQztZ94IkQFm2oUoTS5h0M5bgJmU9LzOeadM+ocXhYI+v6z2eVDAUNOSVu4KGU00VVyE
vTi5/IK8gaJbfgyrWZrAGO6GB7gorL74NriOh3qRMyJpdvXe+yYSXTzt2pgDcX5yEjfLPMRsn5ys
SquPqaTSyT6awZ2AYKFVEfDb64yBbGGwz4yp+Mm/tCWXAlck1kV1I+r0vB0vZRJnIAYervkkRqj0
77nc2L88K36RFYXVKPPtYImVOzalMTJ1GZUirGWhrM2mwtEEqHgsogAS5v+Ctrv9LXVRR1XVUY8B
+57vor3aEZzA2bWIh68huvMMmCntSfFaBQ6QgLPx81Y3nF+/cGd5Q3dGvjhszcQAf/Anw7zreUNs
vrttbkVZG0b274R7A32EZUqdJaw4hUNys358tIBEc/xo83neUpUsK9SxBnYhrwBzIvjYQMGPZlwI
ScNLTRj+6bLtSr8531gXPdbtQcD9W36a2wDd0QlP3xshVx7P0XbFrlqvhBeQXlhSPlWW8IsecNpX
+FmzIBVS2LTp3l/aXYYMzvcNqjQdO++ErLytOuTxt7cVl6lC/e5CpXE1SzmBQO/igZ5zMWpU3K2q
1EArO/PLQW9q84SY1hN/3WHLGy50zNEPJXRDPjMPxBCxLt2uJTe+Jgc32AyQrJ5ybyRRLjOjPrBY
lieG0X8oW97xC2FpZEd6KIfaCvhuAOkjTMh+bhxM8zgg3Byep/txxbRfb/TcLfgQobtMWrWBt4wQ
sCuQbgvBh8aLlp7qFKhzbG6GkhqEzO6zrHarnIloHCUPI/RulNzcE0pwbZ3jDvV+wkmquUx3CRSk
lSfgArb0cfjsNw32+sYePNuNV3MGdOAcfZ7o7PR1pMVeZf2czpNx+ETuJcO7bIkVSXHL7Sd5r60d
mWu2jMntCp0IArENKSA7l3TaxMjo8BH/cek1sjaeQu9EX+Ba628lOMRwx+p49Rcuo9PjCkqtvYvr
x05caemvfCKT0tMNIRGFO0D8/Lk5G6lvIcT8REmgz+s1uGNLimcxGrsXkCzi78fn4Lv37plJekJd
dHjjFzNzz5e1l4elp9cpeufuNA9oTq+sukZywo15S6TtIiqq5tbTLRbvqL3R5D9OYgKzUROKBtfY
SUpmmd7UW78my8CN7LB8mZ/EdpIcFTztrmNf3hzpjqUpGtXTFXRw5zU/35/8UV+Y9i2M6SO9OuIT
04JZ3JJW/54xHbTS5PtM96wLYVND3/IzZW8yOBI7KzCUG6nXnYn3XBlkWb1I0CTE0M3nIpbAChUZ
vk0us59xW72d0zjiaj7UvCiRXXKTo06UYxwOGeGzuZJe/JjzymjrbAZVwaDAsYLrze+cEyFtZ1zg
JhETxasRzxYTzeSfx6zzLL+EgCUKGBa3aJEFTXw/tGD4I3OL25gRp6/oI9RxIN7P1oCAjz5exVsU
bkY+c8RcCyBEhq2j219Zu+TdLpW7jbvfauYucNavC62aCLu6asowMHhFlBN2c1ttQptLOka/wlaN
94idploPKQDGIfEqe5Yr2EsruUsdrHg5Va3xeY8j62c+KwYU0xmiMwHo9Lqdr5BDCDCFGc9DrFZn
59R1AIG8hFTj3AGkEqT6LUa7oMhXNeuLEXx/T4BfKe696TvfUbOTK0e/XMoDyV2/tXyalv50Fb4k
v4JyZmj7bx23eMXM4t6sDT/DqK5ohmim5BSodkBJi9rHC/NTjC9pxURu2AMddoflfKyHQjqp6O/Y
AwmuOhXvIxTDMHlXQOr5zdp8yrRvm7IfJ7UHIlXQtixthtczziqYfa8PeePbE5LzX25uCc8g3uoj
gyTyLwthE0Ztrytz+jUV8OR2EztlPgJAfjA8jxWkQY1//1h97tciupA37tD/o4uluK6q3FAmqbn5
wD6F0iv0P7VnmON4t4Oid60QRVHBRZPiA1yieF8hzDQrBYJ6zGWPVix+SFznx19skVA1amTBriJf
oRl9DG2EuVHwocIB4o7XRWOfND/jO25wv/Q5Uz1oCBzfNuMsongxXl1lFsLBBy5zGfmi6baXjxFu
QokrV9WGlAcP30kPDFL6tlJbr8fzXB7CH0djX/Xqk+/z0iCNem/7+pwkcQwaxhKn9PVcsZ4ykj05
nw2ifdoRnaLLVn1LE66DyvXmXDgU93lMikZ1Fpw+gS82yOzS6tTKezMaeO4bWYUUhMbTWhcO2p2S
PRkOlPG+3UbA4iD0wnh0E1Pj+p+iHVRWG9aIe3ma/JejdIMpNvYkKya7qBcIz+x6ejilnkZqQjT3
cWsphAmVGqih4tA/ae0tQp8DbRNZvHo2ayBtLJLyV1NXB5UTN5HE8Uf+dKjf5w3rzGVnwjkMPPwo
HUpxgLCEW7rVRoGQpCCHoN/O5uHZjDXZDBb8JngviZtYloUKqDHlpMvIBrl/sADt3RG4mhqITwS1
wdUrI/z7CDEUs5uROEDf9lq4HTwEyfZYKM0Nx2rIDTPlzvur7TYecXIib1hlPiISfmfqIdg1ZTqB
0/JXf4bjLJuGLlhv9dK9dWpPU2O5v/3coeVRFPaUJ7xYx9i2z0VIDXagu4KAabCbV86Qe/EdWNdG
Cq9kFf5eoB7Vm7VNGWte7GMOTCbTfO4nyB9e5BOxKsMPFWrQkv+JR30NbOuGQ3WeYSIRkha6geIe
LYfBC0LAW+HtCiVa8+GwlWRd8q3uNg63DWWliZpV8RBOb9EQ01nDUc97bl8x4ctOUiApSK2sw2CI
J6R09gBwmbpKFHIgJ3IFgSBxfNIio+ByBebB2JLXL8sLhePXECxsFnGGsnxkmzNxdHasL05oYUaA
+IGrmEZfumr/ZWfvhp5fLcNZKbbW8lGaZ2TOgF7+p59BfEd0tYpQca8FWdn0HT8tw6/gR8ehk+LV
yw6rQvbR2/LrYAON7n/HR+aJXoF+GshbfIm3ZSeCt4iF57zUsNABnioe2YsSPeyfDy2Rp4wOx8Z2
5Z/eMm5hxIvSWThffqXop+fYQyP3zZ/rwhOkGxxKC9bflwmeeh0/3R6wTSxWOc0FesQGhgr7HMqG
Q3IrbbTTebIoNCoNwWlzyOR705F/xI1AcIKDwwRv5324h1jw8cGG3Fo9L7SYhl0oFfHleZexgv89
926VE9gSJ3Dfkd+o2SMEoc8os+s7VN8r7VSpmSPGD9mXaginLp8N+FVlBb0PkcBLGgnaFe4NOr6C
E0hrhvA0wzXnRTf04xt2f/qxIiRQyCjJ7OmFYARBDeCbb04n9Xs2cLwtFGzcQzoG//jmJm98FRP/
zHde3SeYo0kZM4SFgFCLHnDTPWi0WHilQhBolYL03ZaFa62dRGhuMtHzNPj8MKwXmFoX+KhMmgT7
rfHyJ6dIADJAeEjl+LfWZMHn/2A2oCXWG4qnnj+0CL6lgExEZjtSGUML1reXPlklUfruS8Ag+aJO
VmqO/5F4BjARd+dMROft9dpMnhAS9RXiZ1jIht5CO3Hj7LKnoT0DZQiL35L3BUHnpfRFVmzbwx41
chAURHObKl57IJchlji/jeKfDDKY18U7GTH/J5Q/uqS/6E6PxauyzuPMtczvG3gyLn2kMJYXR9uo
/12X5BCybVl675H3xSvM4LyvCPUjXsXLX1pewxtwU84PtCT0fAVLfKxkUfxy+4nh4f7G56fLfRwc
dcvY/fKr1YEynehVTwq3U+Zs5Gygrm3fBcRYyb637HOj1pcX6lZIS2i0uflWnCqlmv2TLHRkMTXw
uumKeKFx77L9m0PN1g0yZtmUPmIetdnK81K+wfnu44GN6GLnWVeqyb3OagQpH3mWXGdR6H5NOIJp
36mQLPWCr7Gb7FD1PBdD+MkCzjlV2qtnizi8i7ksiJm/GLjw5WBDT9FOMSUxz1EPv4lCHuqY58SP
C8ZCKpI3uMlKR4fUgu6+tWFI6R6DxLqZsLwkpgxH0NvC/PQ5JIvmzXPmoH6ZaK5FBQT9PNTHxnMI
wwPo1ZOJpAodErO8giXW8+S4Wkh9ua7+Ang9xkQ5iUOGDn9lHc0FVwpHzvW7a8MzOR0tCtmrQ7is
lXLdQCWLosuzQ7BzE7AgFye4E6Ffx/TQ2jdf6D3B7zHIvzWCucXc66N7VgNo02o1Z+WxvEc68XNy
cJIx2g0/jx4pTWNj/s/YD5H2uWXFpsOxR8upiCwwuSQM4ZiMdidbnUziD81/C8YnxLaCQOW8RsSp
rMABo8AbwFTSfj79oGMYUgrbQu366ACv0SvByeAgXxmU8a3fzcrI1YoWqpy/sNOIHYUhV64m3ynn
A1fUBLV5xb/HZCI06u5aHn0oOMdlh7wLGmeJZw1tcQnIbCZ6tEWIjGP1CKYOB9RebHncikNWMlU7
NA5VP79LOSPnvUgRytIG39c9gdLC2mu8h9m+0KrgJMZf6cZMMrPov3ee936a4UHVHfWhDy7qWI2T
CBysNys6lW24EAAwlhO4cOLM0GGofEHarhfrYgWneEpiUm0RPC5yWq779tPJW9FwYPQf6HSKTO0u
0DhDr5CJ3MSffAr6DZ14ECOfbdSv/+Lwkd4K7AJy486FcWUjWE6cWOp3vlUGIuh1pNJUjc/d1v+j
C/giDCU5MI3dGF5AJCDLPBftjAHk7FFwUXKZR1mTZ6vazjHGaemFjGjMClkdQzmEfdyI+YfLX2K/
7p5LwXRZyL4+ms2IX6iz9XJDC1EwPu0dBH8paR3CjM/0tIW3Ao1Kiotb44z/F/NlMmRu5zTLCmTZ
2HH7NLjY07sqKprQUt42DlPnTpPI6TupdXSlueySoR2i8lFSXcpU1StvVHSX6eYuSU2K0UpbCon5
ifog9nW1BI4yvGc6MpbSft9qtz3tYtuMFyoSWYhShz42udXBaJPqC1DJWDhGqe/pVTML9GlySAQO
4XQ6+O4oQQi8DxlaXtYF75r/EMVNSMtw9oDJTpHGy9bJY91PMd1vcZCexslSziIJ81s5Ka91691N
fxrc2g52AYvrgqRCnTX9Gpr/y1JIWRikOuQDrrBjLhOnk3fkOIBYZ/2Cis6MjkJoh+XGUWfjCo1d
owWYNL5L3WxvbCnQETu9M3F0XisgTiqrgzEo7md6qYnLN1R0NwQ2yz7AUQ2OxGtpwHeBnYEIUY81
g2VYpdGoSNa2C1yd2MniYib2hW7evp7hFV+7QCiBf/r5NRE+PPz238wgrze+RDdHLwBsqnglBC6H
v2s7lLKPOdJnf/j3B+cXv3rEmjmNCmMjnwDAu93cqRtZX94vrwGHIMkm3rD5Om1PYQ4lHYpQEwNd
SqLbsrf13lf7jLqAwEZf/syvhW6rT6tixYl9oECYchbLbfzSDz7+oFBlbsKbMQLMJgwwUIrKJK2i
iPgWpzAYqvgUipH7snwaiXmZ9JGINXhIJBMWAqvZO1sicgJ35mqUygedPlaPvuBLRasFGoTJDFpz
bzEG4nYQ9obIFTu8iXdw6j1PcN3bwW9uqCo3pSp9pMP97DSUyC+OLpe7KP2WqoTvBygrQfpYRbuH
EPx4ytG+pR4WGIKuZQVmGryHOmuASmoBhZ01EQZrNWbhPgdALr0ysOHKDqtusUZOqDw0SVph/abY
yOu4iO3oAG0JieZpi4WYn+pPizYbNqsxRAjcJllEbHPpLuOrZStgN6g9vMIJqCUIv6YfV/zeVWJv
YX2+zc3Irfc3URhr9atyWqTHJ+ci8PQVJlY9GHwUWv5RIrUuZE5bntYVOTy2z6NoY9q8/sXhZ5W4
5XB620kwC7mSaK30yApZ+7IbAc/4d9AgwvXZL3uoR7p5kyY7h7RgWGSUpOSrLBf1cfNOrn6NwGee
xP92LxtRLraWmnlWl/KqLSZBjYL23xtmyDT2KaYdv0CD7QqCOipc0JTNsRF4bhj2dci3niLMtfFe
eE+d6CYVtOxR4HUGvtXgPbNN064Tl+5GBPUYL7Wdrbc2XMOYsy9pk357fNJ/c9X3Vun+zsVZqGIx
lY7XFXXxvgk0uTV5pRMrpYpWP1onUlvUSgj9cUixAThVy8w7dpZEbesHZze/VcO3soWJRlYUeHHC
qm5T0ATlcN0tlZNt49NKjuHq550vcAWpSUjiOUJcfiVk+aGsMG7RizjRCY93x65hLqTkWktmao2V
EGG3pDbJCHP4WeJjyQ2tHStw9rTkYOyGp+vUaZaIWVAjCQISLDqmrilb7dbp0vIKdZQeNhH4DifO
3wdKeVDvJMQ3rtKjdGDuGPQFRG//SZrZkhxtk2YHmt9T8MXeEHnW2E+67cB39DG8IDyEkvkXK/x5
3eVVrSVFOVlylv2pHgioO543/9cDuJMd14wlCHcfINOXsSxxDzSBdrX/ERPKjrpJMwdIpWRDmBB9
IH26atMFnf+US1d97urRtzSAR1ejSwGWr+JrNrbIploHAVdqi2Kl1wEI4kTp94pnFNDjivUZenQA
8OjcZmaXRhfoJH3CkDClTDgncLUbHIAnPYsHMR+MuU7kgEqbkuDpMk/HyjBf3A+oV5cRybC9UdND
V0pbmA3W642QOnZy2rYauf7rUIOMFRiYtuq7d1qIWwJqZyqUaTlsuLyiIZSRY0/EqNuUXkfvdKuv
xkI/+mELo4f0RJME5WxcsRFnEcz6jzQzXWiGr+HNqRVZXQeOOZh62B6XnDQyMLsRGPiZoHDepakh
ny+b8Ukc3/F6ye9QDJBtwmh7TrR7f2wdEKV2gEEI7Sjku17PLNXmE1YR4JuN2OXEVhofAeL6Hhb0
WN7PQET6wlH10ePb73nWNTK2Uf6Be4jJNsw4z6CiKTIQC//G8YTd8oQDXvvCkr6GIDHsqT/MHM5I
mhbUApJa1U+HlrvHbO2CNFTOQOyMHC4A0gAZKQIV9yaKD/U4Th0DJoShOZKiONqsw+nwUAiFFxq6
4hy1fkJVoBErTo0SvpT5e0OD98Zy0FRZRXeFfGEbO+t+GRwsti9Kp5xRGZGpXzRtxr5Xql6wP3gF
y86E59WiGTX/rifCplZKn07QdAdrevjZNq9WZCnGTebvq1UcUH8D6lfwHgzoDHoRkO+9XEae28vh
yRhHmIH0DnokvLp0kV4djM7LTKBnjgZBKnOo6FEE1M0pMWs/sHeUtS1Wt60zcyGcnSYL6wCSsHho
a2QS8wAp/qabDiQsauKpJEst+GiFqZrDl+QLg+Rh3/CjY2IUHkV9grAj3Pm9flmABnpPc7ilJAmP
x5e25tUYnughrkENEPP5D9M+HMAWj+pqmVUa+xrcGnrkdHa9/yJeEzesJf+jGjQc7MCb4bB2gjST
o4DdCOKMyI+fdXkigoAlHIDX5o3MFf+CgJXXPgkRJjSIblas3B/gBC1vetEgL8U6wbJ0dMu1iLZG
pmsXKtnneQFUfzUgYJBjU7xhOKkyTw29allMp/M9F8GLvYLCBcpB9NIQHY540R2UEd5zBswfzcmB
u3idc0HHl6H2Q2u+rqwfdYkNLXQVCLnWbUx5F0Sva8IJGtIs3E9wPSDbLZR9DLsm2Bn8aJZtdczI
NT/lJJvjHryFdzVQoUuGn8m/ws+BYRhEBOyRFmRkEld9JhIj1Z8qS01dkrhyX7zRMcxwT30/yRRe
tzRnrREXRQcQz1v78D1K8wbOCfyh9BT4PrJ6xkI0XqwxmwVHCaSGkoNyb6PhgtcLV1Jbm5bUqELN
vPWgSuWbS+GwcxXzLcMj9HGzW6cQ1uhKqDNEIRHf4+ixHTXJMeB45EahtAnsCc58OBAQX6Ds308g
fxu0T4+swOIUmP66uy9/WBPPXzGONC6Iny3au4KPvwmDR0kVIs+dv2F6ziTC+BlhaBAD1zdHGn91
BZtCo+seaytpmymRS4KsRXiLYuVRoHN/j7shr3w3JHDbsWj6dcBpa0CcFrIojMjYFh+UBFe0WJS5
M5O0V17zBc1TtgVmtBbzhfh8rDFMrYH5vdF6Jh/wzP7GFKN4FSXYf6eLRq2vJYGmlNbeBmYgSwYY
D5gNCfFxzFZXaVapgSw+vLY4ybYqkKpc74XPuSsfzGmzHLHNXO0d0hn75td602B0VvoJaJbURrFO
a1VsbdPQnzFapivDjjTOH0EpPfg6L19Ipq9vg+81URKKixbq9YPTKS1CfIZnvRv6igRmNYDAjG3c
RxgrEFdW4xF9/YzbczYG+w56CrPWerxWwfIKhiwmSVkZklfepB6v3WnzdZgdkp5b8UDhBPEVJzEz
Q8J0u+i6G3Rcv3tMfAeabGV9+dJVHwWlCqX249A5XxOWswH7Sa8ansBKhz+2kWre8e6j2bppv5sd
SvCmF27L89cp4SIVS4vI/gSgS7+b8n1Yexkrt1aUK/wRf2bGOIk/3BWyVNAXqlUCBqIdq4Iuf6Qn
Bd0EESjRioHHlMS/n72z44kz+/Y++DCd4wL0NLBEkJg/Q9g7nObMWkXJ3bnl63umBhgn7JuVy4eH
206+r9c76JqVP0Q/3k7ddXroMZ2jlvlYw45H9mo1DoDEED/whtO8VJRBtSHHU9cAkOOiMd1LC/l9
3E2efLwnDILEZY9o/rw/TUxyj290fnZiF1YQd4aEaZc0qDJuzIzNdxWdPc/yI6no6/+9PaMrQO7k
5zQ6zkTuRoiTS7fgM2/Uqe+EKVK43P6prfdcxlvRHdsJ6wFIi7M/6Xt0QB3HyuOwYle+g7ibuAlS
YCgN49q01SToNKR9YcQUD00jSpUxS4WZVJ8V5CE8TXVwwAL+ej6ESUK7+iVI5SYUjGhf7d7dnlSA
B0HncQILZKDJFR24lENbnfTWVyzNYT4t9yLXYUd4zpxD59nypMf+BOoi2/8WI4Qdbn120igrQnLn
GSrZAmKFINFqY8CJ4HbB9Wb7r2H0h+Cdqh0003q21Pfnu9dA7HDiA9uVpfZLpuIW+0a8yuJhO0s/
+MztjEKv19P0cvJRWX3huj+WX6T6CoqNPvMwDw+5prOBiMxkjUvEK0jOVVgVH2vpSjd9mSRK8IMr
ipIACpqdKti72x+lORQJdWdX9TldBzPiW8mgRkaKhwnsdw9/dK5RkJaXc5ydZYj3y49Dp6XDBgIm
gNwMbgEj/g2Mxr/XiER8degn5talbRbneG7AE0dSP9Tn4ZdquEFVfybX4xZPURnc2tLxfQBaqc6w
2h3cwON8AlGT0Mith0oK/R3/suR4k+CFBGjPK7EF1ixvLUwPu36YNDnJ0AYFNJePzglGBrXKAUfA
U+tX058vr3Vg4suNhGNQBHJ5Cc87KvzmzWw2lviFeju5pl8gF04K9S8IOpQMzgIIfCrhAObctOiH
3JR/+AL6wVYo759jkO7RhGfHiXA3lpcKlaX38Rapdafd96w/Q2lu5e1tVqy0B1gBeuiEyz6cfF98
rhFTUdyuQBqMI93lLjSyox9Lwtc2yt0MXyI/WDDRoNVXPMD7k2riKd5Bvm/xSCQ295BgYSyq/tfD
gRzhQ6lsNyDnXKEbh4b7tdfy1eINvFssQLn94LNm64+RwBT8kNMPuDPLbHuqdHNeCh3TpPJ5UWVm
bxriI9C7oODSsLTsPRJtnGKL5y7GYcWezzVsRnq1AC5VMB+43hennAOgge0HVhywrWI8VcFY8Aeg
OCurrAyHPuzdAG68voRnamH7p4yP6hvfbk1eUXx5N7W7+s5KWQ1eWyYfwO2aDipLGfD8qRPg2S7O
OVXfXHQerT1j7rp7x4s7ywskwKTWDSE36yYF/efghIAqJQ44T4L89aGI7H7GTOT/vzUvUIM81ZbJ
u2P8Il8X4c72r0xRdXkfMWUFQsnkPwDdmToUVynUQ+mYaMUVUYh6fLHEDfuNjH41dE96f4mEmd9K
QPmBdyb9mAkXw9NzKVa1Hg1/d/xfhfe1X+F7HC1U1z0gPdVooIqR6ALq81hbw+3mhIKVL2DuPhqD
Lt4S0G3xZNNWGgeJld5PVJO4/ahWEoHKA+APqoR+1IbT4MFCUfn5kpJTykGZM8auzypA4crbKfYj
sjtrmKgL5dUCkVZqhc5jzAIjcPH24G0HYW7zdhuvM7Zh8zh1NLFt7mAF8hz+Zx+cErUnQCOOxAQW
dBxUbaF5blRgYGm+YVf8T0TVJ8EB3LWT33fzgaMWLO6IRZk8lyETU7x5X5z9BbEyoY2/RaI5aP2e
pbmBaOoT+05EBX7UwD0LsWjxPMx7IQtp2bksHb7L7iR+P81wVTUYrFRfYYXd8ONOX6douKvYFaNm
HGyVOJ8v6Mol4W2UktvQv1p+Hq8O0X34pFvqGe0yGyt4yek/LKHv8VMnkD4K7WoZ8iIZ9pY2db5E
LOwrxeG83n6icNxZA7UTTAy66+h1FoFEbykYvJySu/l0AyMaMIsUmPuwG/L1a2M1H6LQvqmmg6Bg
7cAqCC4uCySwatR9JH9zVkKGHLr8o1E9QPfIVdVJAT3awIIi0UX9ZIep2BhdU3hrOkYTUEBBUSqn
j99ZQ/uOr4IBBtYEGTWXVMbm+4BHC/Php7I4E4erf+NUDtZNxGe+eudJKlInQo4IDnjd9ccflOmW
SIc4ai0qwOZrcC3chMNtJ5PvEhXEMEfAEL3ngv7V1FrFCBpG18N+ht6jkg9D/oIPXaNCA5ZsJPr/
2dsTCSU5KJ7Z7wmdbNnY/uR8WBR5ksDGw9wS7SMwyLDaHABmm/tFFzQOq4WRstB9wTIv5Ge4Gdz5
Zy61CU56r33oZpVYOV4OwV0fUaZv7qEl2RZzUq0jI3k5CFZYJaCjVGq93dzcBcinkoGZASDAqSxa
zvnWQFk0aoWJS8O5PUAS7gZeJY90T/8Gm5erAByco56ZC3gUHRdhb8yy0etEEBrbBhCg5Vs6H23H
z65K3dPW0HU7GRt3u1mJ+LhXqfai9BT/mGCK4FfI63Am1O/Kg5ms5ZY0h94t7xhYzCaPNk2WfTJh
wzpBGi3z4DCu4a5j0HAOxSrxGTeBrHmeMNmqdh1xcqEN4rjnL+NzQM0axPWGd7vf7XBsKEZr6ASz
WvcoCW15TO5pcSj1dBzBmuVsfu+faajrowAOy/WjxxUJb2VEyg4PkN+uUZ6A2ZfhxfBghjYU2NbE
efUcEtrEVuNmNptUwuy8JHxR93lm3i5BJvJo1SgbbV6Jt22WkKb9ZEWx4wHmyQMKC5pSZopr/DJK
R2ABQKl+OUjrK8k0OKqE2vlU9OU+jde+E2CkCVxvv854N9KPytXRMiEkty9a1ZaSR/z+NhCpQ3q4
XHLByNlM6yiyT9WRoedLQ5uxi4Jtsgz7M3tGpIqOYNAVCZr64LyL858bJaq1BhkqlwBc0jfmzoqe
0T0xTO00Eq4UfFVs+vX2ipb16LQYJXiJQhMPGkmdFSkWB4MEBAVyz57kBEUCpalbfBQJkHExG3RG
r03LZ8L4lhkwCBHG71QG1n7SXbPS8nBpD6eozQPsJkEvoaYsIswYhRHRp3pITFN0RHXFOpUQ3Loq
E5Ihcwyf9M0aUFOO1dZGC6CJm1rQzwUXWuJf21o9fGtucvD1KX1WByY/Hq7Oi9szOWOgLKJw+HvG
wINuzYHnaieJ2b9ryTx3A2D+JZMDww4TIFEslaqEQNvTkg+Gc6f6pwCUAqbeYkXyD0xwBwdMqRDL
oNdXU4wFGhLWap9qH8AYUfUGhNYdiigdk7SP+uG7lRoXf13jP8CbwHYbqAnZHuVb0sBkCaCFs7fE
hngp9kUeuJO4pt30l6rQMfBNPYIFdHkBtFZ+Kyq3aAjOw/vgSYhDTZCYPAq+p3Qj/GwavEdhDzf6
bknw7f2Ns4elE2szzfn51JxPuIT2syardPVYGvaiRwamdlAhz8JBFF2XP+LJvtV7abXQbJqDHepy
gHx1o+gmQYCEv6Oer4V/SJ0ejlb/vWVw4dyjS2k+qNa1vKRK9XsbcFx2YVODjEgCp8hKPz5PRSKf
4xDnYieXEqu5hQPpXQ8fEgiwHMX/XVjtJjU+3H8Att7pFT3yGJIgQWZPTU2r3FPTwtSNUw7lKrdV
DxAa/0Epxn6GWgPcyFC9RinqaQbwMbjb5QfzfCZ9MBTujyuzqx9tiyhkBmYiQv+Mj8b59kyuWZf8
3qdjUlpe+uDy19qqsrHXU3BJvB1pI6Z+MqbMgn3keAreE8hR81rMOahXuFx4aymGp/1kNxRC01Y6
zBWk7fwkuJyg7IL2vrXZtnmhMoRSe8/sZPoGFLooJ0ioD97BNymejWd9bnjZd80mNfomrQvBFadW
4SapoMh+Y/Qw9VPAhsVtQKWbT6awKukRsWyv8hKhfmRCQAtCVUBqY8rQMWN1qXZG9dLNKMZeGrlr
H8QwMMVul8Q0DBroyi1SSXL0o8BZGo2AHLpxt1rqOGuD60WcY//WSLeYI4WkSaR6+SWMB0I6vNOF
NEosPEOW5NZDkrveVIE0L98/aX9n9Vv4R02jWNq1bFGBVD8AE50yMWm03dAJE+RqnLhO781qXI34
WtdG8jJY0rC6TKJAwbTc8T7s0ZZLgPC+8grOKfBpHoHiWWji4dCLO8Hd5fmC1hIoaAkk08tdXZdH
NsU5/94S/AM50YkTenQm59gZyQdjwY+eDBgcPhBaXi5boo4bdlvL9on24bUsEaGdK8ITaxJXeEY2
SQmiQZqzbDcuplkjbYWDg2PFB/8yf3ThxXJdihRba4Aa4af3k0VwkRuCMPPv6yexwGPEzySb66qv
xBp0srvSRC2PikBsDEURCiMX3+x+t5gYKj/3ven/moStExUpYRW0c6mU8zmuUqDs3sR3hlMuSNHj
movCGacCy0F8u/rS76YOafYyTCj4xETaUbOMXtaRftSKr2Qrkw+j5dquww5ZIVuFN8FwJwWHy0AJ
oFDLyAXgsS4tDAIgI3/BMCKmIM2E3xOUNa9ey73ZfU0wcJYnFHiabk+Fcum4bXaGTiU6Sf2biohT
VLv8OBqGWLaPJDGGlW6+5Yu6QvH+nhkB7TsWN7XJUsiz52b9aq5e56pnoMu6TxxjPWbOSFcDPpTZ
LX5XZMlD60U0vZwdBjF610tQba6ywEC9v27Witf7i4mC6UhqzKQnRlYpHibJRFM6f0oBwo+OweC1
Yupl9vRdbyFbx73x+L5D+MI90KIRl7vnqGI/gR1HSg6lUcU6Nh8jgt64DYE/Vdfhhhdk4firXBRV
lfGw1vfH6WbxgneMoESe+hC371U4r7wjDgzuofjJGdveDOJHDsgABsT4GoWBNQWB4v/1AFq1nQ4W
ojRhNU4dS6md5GyygJHIEAgOqjenTkRh+yVJeadHFtmBcMJ7+3e1a9pntmebcvrJFnFYSZfhgUZ5
ZGgVBg+TOJQOQhUfYUaLPuZIriK9cusyZL3cViQgUj8tQW0zSBduZk+EHC4nNTG78NTo9KNOb+Ju
1W9pVYfpdwgrjMi3+nrwZcKBHNqria0NN7QOx3MADJJ7CKxKF9odVDpigha1iyOadnPuCAJn48ED
NqrcNNzCoAwfy6NgKie+I9vHMt3b2zQxUMtj5ehsX1ogPBJRS8vs4Duxq+Sj3YfQo0Yw5MTTBWFa
O0oAz2YM9UqVwMUgkx1fv+vID1vvOY1CPQ75eAM0loVA0Zyu/s0hd/PqrR3MKr6hL2ZUI8YD897v
tTIF9l8UVtpENQtQOlRrCOtlpvKRuMLoeAuYnUX2a+mRYV75f7RV3RKLUhIyz+6HiwAFknUdMsdV
v0eUV0n8aUc4Wh3We4kqitmcizKhcquJQ0oiPGm7SdGQeZaFduy5c+BHgAHTt0FhYdaWiPwO5OD/
e9DrKSeieYji8FGhQPhjW+Acup0PsdYUMow+Y53EasXZF1Re1wb0JkntOgu3K8kGRdNVONpIwuIC
i30rWEbGj10l7H4HI3dlnQ6x4HioECs39bJtIw4Jj5X7dx5LzeCzI5SrTD2mFZSRbzQ6KgIs0Jk7
wl3JPr6u3fj/pLalk1l5mwG46b4+dnCAIdeGStV3rjc4cQ8lW7vyBGCgAVXCnYGnfIarWluFj+is
br2AT+7d51yTbKnSBEe1PorYXip19gbvdPmX9HcoXuTPThquW4rcMwQFGCWv2oQ+EYxLfAPNtqgi
MoYb5apFvM+4E3bLudk/38lcLprRKJRYcoUmeOHw+sX+M6Be5qn9YbfuR3VBO1IiXhfJ/pKfOLC0
46+kF7C2bWGQ8OaeGMvcP0O+XioFYf/uiBWFf77YsjKNgqC+XGGQcAJaA/uDfvThG9LWlVwcnOI0
e8DS0lEfJF/QtnYnJ9FkPdbtlTRIl7PVM/vt++zUfauRZ4kUb6MLH71Bu2c+hwiq7AM/zOH/Epqg
lRMvtfF2WiOsmZ/BYf1jZ3h7SVsFhFDYeY6cb5D3YfEmJz2anpPFuSJHfefOqqJCujbx3r0174LU
aUTfFs/l6beTUw9OpaVG5azY0DXN+SQy9OA4dkFjpt9gmRJ1GidIyUFd400aIdW+za0o0XlMlc+z
dOoZxtA8hIwurM2j9Ct/f35NWLfMF3ONlsfnrZlnj8f0OWaQiJxaYeEYGYHmDF8Q7b5PfDnHbzQX
1iL5P5/PNUT8q6UORGABPH7lw/SfptkLbII5a0snCY0ceBXZcA37JXvCtx+k34lkUPLVgzD/VzLs
7583fWvJTz3uiRp52tOtSOL99Qz7E2Ztk+Q85UX+mwQ5dv2csq0qIB++uS9LNTsrryzrFSmO5Esm
gHn8QZAecQUvUVbixEKrfNBzxPLwaw7glu5zcQLl7EY7ayw8VrGHHmgT3mwl2kPz+9HIXftiCZuV
gEP9tgDVouhm92oK5D4l+2x5nKZzotor9PJnUw==
`protect end_protected
