library verilog;
use verilog.vl_types.all;
entity expand_task_vlg_sample_tst is
    port(
        clk_50mhz       : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end expand_task_vlg_sample_tst;
