library verilog;
use verilog.vl_types.all;
entity mips_tb is
end mips_tb;
