library verilog;
use verilog.vl_types.all;
entity led_vlg_vec_tst is
end led_vlg_vec_tst;
