library verilog;
use verilog.vl_types.all;
entity test_OPD is
end test_OPD;
