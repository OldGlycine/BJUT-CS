library verilog;
use verilog.vl_types.all;
entity test_timer is
end test_timer;
