library verilog;
use verilog.vl_types.all;
entity addr_38_vlg_vec_tst is
end addr_38_vlg_vec_tst;
