library verilog;
use verilog.vl_types.all;
entity controller_tb is
end controller_tb;
