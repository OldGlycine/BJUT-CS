module timer();
